library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"AF",X"32",X"01",X"68",X"C3",X"D1",X"00",X"FF",X"77",X"3C",X"23",X"77",X"3C",X"19",X"C9",X"FF",
		X"77",X"23",X"10",X"FC",X"C9",X"FF",X"FF",X"FF",X"77",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"C9",
		X"85",X"6F",X"3E",X"00",X"8C",X"67",X"7E",X"C9",X"87",X"E1",X"5F",X"16",X"00",X"19",X"5E",X"23",
		X"56",X"EB",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"E5",X"26",X"40",X"3A",X"A0",X"40",X"6F",X"CB",
		X"7E",X"28",X"0E",X"72",X"2C",X"73",X"2C",X"7D",X"FE",X"C0",X"30",X"02",X"3E",X"C0",X"32",X"A0",
		X"40",X"E1",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"43",X"0D",X"BC",X"4A",X"6E",X"40",X"40",X"53",X"54",
		X"45",X"52",X"4E",X"40",X"40",X"31",X"39",X"38",X"31",X"3F",X"BC",X"4A",X"6E",X"40",X"4B",X"4F",
		X"4E",X"41",X"4D",X"49",X"40",X"40",X"31",X"39",X"38",X"31",X"3F",X"54",X"4B",X"40",X"4F",X"55",
		X"52",X"40",X"53",X"43",X"52",X"41",X"4D",X"42",X"4C",X"45",X"40",X"53",X"59",X"53",X"54",X"45",
		X"4D",X"40",X"02",X"3F",X"D5",X"4A",X"32",X"40",X"43",X"4F",X"49",X"4E",X"53",X"40",X"31",X"40",
		X"50",X"4C",X"41",X"59",X"3F",X"D5",X"4A",X"33",X"40",X"43",X"4F",X"49",X"4E",X"53",X"40",X"31",
		X"40",X"50",X"4C",X"41",X"59",X"3F",X"AF",X"01",X"02",X"04",X"32",X"02",X"82",X"81",X"10",X"FA",
		X"C9",X"3E",X"9B",X"32",X"03",X"81",X"3E",X"88",X"32",X"03",X"82",X"31",X"00",X"48",X"CD",X"C6",
		X"00",X"3A",X"02",X"81",X"17",X"38",X"F7",X"21",X"00",X"40",X"01",X"00",X"08",X"71",X"2C",X"20",
		X"FC",X"78",X"17",X"32",X"02",X"82",X"24",X"10",X"F4",X"3E",X"08",X"32",X"42",X"42",X"32",X"01",
		X"82",X"31",X"00",X"48",X"21",X"C0",X"40",X"06",X"40",X"3E",X"FF",X"D7",X"21",X"43",X"42",X"06",
		X"1C",X"D7",X"21",X"43",X"43",X"22",X"40",X"42",X"3A",X"00",X"70",X"AF",X"32",X"01",X"68",X"32",
		X"05",X"70",X"32",X"06",X"68",X"32",X"07",X"68",X"32",X"02",X"82",X"21",X"C0",X"C0",X"22",X"A0",
		X"40",X"3C",X"32",X"04",X"68",X"21",X"00",X"48",X"22",X"0B",X"40",X"3E",X"20",X"32",X"08",X"40",
		X"3E",X"10",X"32",X"17",X"40",X"3A",X"02",X"81",X"0F",X"47",X"E6",X"03",X"32",X"00",X"40",X"78",
		X"0F",X"0F",X"E6",X"01",X"32",X"0F",X"40",X"3A",X"01",X"81",X"E6",X"03",X"FE",X"03",X"28",X"07",
		X"C6",X"03",X"32",X"07",X"40",X"18",X"05",X"3E",X"FF",X"32",X"07",X"40",X"CD",X"8E",X"30",X"AF",
		X"3D",X"20",X"FD",X"CD",X"9D",X"30",X"06",X"04",X"D9",X"CD",X"C6",X"00",X"D9",X"10",X"F9",X"3E",
		X"28",X"07",X"C6",X"32",X"67",X"E6",X"0F",X"6F",X"C6",X"63",X"77",X"01",X"02",X"0B",X"1E",X"09",
		X"4F",X"57",X"70",X"06",X"03",X"DD",X"4E",X"03",X"10",X"FB",X"77",X"59",X"06",X"FA",X"80",X"77",
		X"0E",X"10",X"06",X"20",X"81",X"80",X"7E",X"FE",X"6F",X"C0",X"31",X"00",X"48",X"CD",X"C6",X"00",
		X"3A",X"02",X"81",X"17",X"30",X"F7",X"21",X"00",X"50",X"01",X"00",X"01",X"16",X"00",X"72",X"23",
		X"0B",X"78",X"B1",X"20",X"F9",X"16",X"3F",X"21",X"00",X"48",X"01",X"00",X"08",X"72",X"3A",X"00",
		X"70",X"23",X"0B",X"78",X"B1",X"20",X"F6",X"CD",X"03",X"02",X"30",X"22",X"CD",X"03",X"02",X"30",
		X"1D",X"3E",X"01",X"32",X"01",X"68",X"21",X"00",X"42",X"06",X"0A",X"36",X"00",X"2C",X"36",X"00",
		X"2C",X"36",X"01",X"2C",X"10",X"F5",X"21",X"AA",X"40",X"36",X"01",X"C3",X"17",X"02",X"3A",X"00",
		X"70",X"18",X"FB",X"0B",X"3A",X"00",X"70",X"3A",X"01",X"81",X"07",X"D0",X"78",X"B1",X"20",X"F3",
		X"3A",X"02",X"81",X"07",X"D0",X"37",X"C9",X"26",X"40",X"3A",X"A1",X"40",X"6F",X"7E",X"87",X"30",
		X"05",X"CD",X"5A",X"02",X"18",X"F1",X"E6",X"0F",X"4F",X"06",X"00",X"36",X"FF",X"23",X"5E",X"36",
		X"FF",X"2C",X"7D",X"FE",X"C0",X"30",X"02",X"3E",X"C0",X"32",X"A1",X"40",X"7B",X"21",X"4A",X"02",
		X"09",X"5E",X"23",X"56",X"21",X"17",X"02",X"E5",X"EB",X"E9",X"C0",X"02",X"C1",X"02",X"C2",X"02",
		X"20",X"03",X"B6",X"03",X"D2",X"03",X"19",X"04",X"DE",X"06",X"3A",X"5F",X"42",X"47",X"E6",X"0F",
		X"CA",X"79",X"02",X"21",X"19",X"40",X"CB",X"46",X"C8",X"E6",X"03",X"CA",X"0C",X"0C",X"3D",X"CA",
		X"D7",X"0B",X"3D",X"CA",X"1C",X"0B",X"C3",X"D7",X"0B",X"11",X"E0",X"FF",X"21",X"E0",X"48",X"3A",
		X"0E",X"40",X"A7",X"28",X"22",X"36",X"02",X"CD",X"B1",X"02",X"21",X"40",X"4B",X"CD",X"AF",X"02",
		X"3A",X"0D",X"40",X"A7",X"21",X"40",X"4B",X"28",X"03",X"21",X"E0",X"48",X"CB",X"60",X"C8",X"3A",
		X"06",X"40",X"0F",X"D0",X"C3",X"B8",X"02",X"21",X"E0",X"48",X"CD",X"B8",X"02",X"18",X"DB",X"36",
		X"01",X"19",X"36",X"25",X"19",X"36",X"20",X"C9",X"3E",X"10",X"77",X"19",X"77",X"19",X"77",X"C9",
		X"C9",X"C9",X"3E",X"1A",X"06",X"0B",X"F5",X"C5",X"CD",X"19",X"04",X"C1",X"F1",X"3C",X"10",X"F6",
		X"21",X"87",X"49",X"11",X"20",X"00",X"06",X"0A",X"DD",X"21",X"00",X"42",X"DD",X"7E",X"00",X"4F",
		X"E6",X"0F",X"77",X"19",X"79",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"77",X"19",X"DD",X"23",X"DD",
		X"7E",X"00",X"4F",X"E6",X"0F",X"77",X"19",X"79",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"77",X"19",
		X"DD",X"23",X"DD",X"7E",X"00",X"4F",X"E6",X"0F",X"77",X"19",X"79",X"0F",X"0F",X"0F",X"0F",X"E6",
		X"0F",X"28",X"01",X"77",X"11",X"62",X"FF",X"19",X"11",X"20",X"00",X"DD",X"23",X"10",X"BD",X"C9",
		X"4F",X"3A",X"06",X"40",X"0F",X"D0",X"79",X"A7",X"28",X"48",X"4F",X"CD",X"7D",X"03",X"87",X"81",
		X"4F",X"06",X"00",X"21",X"8C",X"03",X"09",X"A7",X"06",X"03",X"1A",X"8E",X"27",X"12",X"13",X"23",
		X"10",X"F8",X"D5",X"3A",X"0D",X"40",X"0F",X"30",X"02",X"3E",X"01",X"CD",X"D2",X"03",X"D1",X"1B",
		X"21",X"AA",X"40",X"06",X"03",X"1A",X"BE",X"D8",X"20",X"05",X"1B",X"2B",X"10",X"F7",X"C9",X"CD",
		X"7D",X"03",X"21",X"A8",X"40",X"06",X"03",X"1A",X"77",X"13",X"23",X"10",X"FA",X"3E",X"02",X"C3",
		X"D2",X"03",X"CD",X"7D",X"03",X"21",X"AB",X"40",X"A7",X"06",X"03",X"18",X"BD",X"F5",X"3A",X"0D",
		X"40",X"11",X"A2",X"40",X"0F",X"30",X"03",X"11",X"A5",X"40",X"F1",X"C9",X"00",X"00",X"00",X"50",
		X"00",X"00",X"00",X"01",X"00",X"50",X"01",X"00",X"80",X"00",X"00",X"00",X"01",X"00",X"00",X"02",
		X"00",X"00",X"03",X"00",X"00",X"01",X"00",X"00",X"02",X"00",X"80",X"00",X"00",X"00",X"02",X"00",
		X"10",X"00",X"00",X"00",X"08",X"00",X"F5",X"21",X"A2",X"40",X"A7",X"28",X"09",X"21",X"A5",X"40",
		X"3D",X"28",X"03",X"21",X"A8",X"40",X"36",X"00",X"23",X"36",X"00",X"23",X"36",X"00",X"F1",X"C3",
		X"D2",X"03",X"21",X"A4",X"40",X"DD",X"21",X"81",X"4B",X"A7",X"28",X"11",X"21",X"A7",X"40",X"DD",
		X"21",X"21",X"49",X"3D",X"28",X"07",X"21",X"AA",X"40",X"DD",X"21",X"41",X"4A",X"11",X"E0",X"FF",
		X"06",X"03",X"0E",X"04",X"7E",X"0F",X"0F",X"0F",X"0F",X"CD",X"04",X"04",X"7E",X"CD",X"04",X"04",
		X"2B",X"10",X"F1",X"C9",X"E6",X"0F",X"28",X"08",X"0E",X"00",X"DD",X"77",X"00",X"DD",X"19",X"C9",
		X"79",X"A7",X"28",X"F6",X"3E",X"10",X"0D",X"18",X"F1",X"87",X"F5",X"21",X"86",X"04",X"E6",X"7F",
		X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"EB",X"5E",X"23",X"56",X"23",X"EB",X"01",X"E0",X"FF",
		X"F1",X"38",X"0E",X"FA",X"4B",X"04",X"1A",X"FE",X"3F",X"C8",X"D6",X"30",X"77",X"13",X"09",X"18",
		X"F5",X"1A",X"FE",X"3F",X"C8",X"36",X"10",X"13",X"09",X"18",X"F6",X"22",X"B5",X"40",X"ED",X"53",
		X"B3",X"40",X"EB",X"7B",X"E6",X"1F",X"47",X"87",X"C6",X"20",X"6F",X"26",X"40",X"22",X"B1",X"40",
		X"CB",X"3B",X"CB",X"3B",X"7A",X"E6",X"03",X"0F",X"0F",X"B3",X"E6",X"F8",X"4F",X"21",X"00",X"48",
		X"78",X"85",X"6F",X"11",X"20",X"00",X"43",X"36",X"10",X"19",X"10",X"FB",X"2A",X"B1",X"40",X"71",
		X"3E",X"01",X"32",X"B0",X"40",X"C9",X"D0",X"04",X"DD",X"04",X"F1",X"04",X"FE",X"04",X"0B",X"05",
		X"18",X"05",X"27",X"05",X"40",X"05",X"47",X"05",X"59",X"05",X"75",X"05",X"91",X"05",X"98",X"05",
		X"A7",X"05",X"69",X"00",X"69",X"00",X"7A",X"00",X"7A",X"00",X"8B",X"00",X"A4",X"00",X"B5",X"00",
		X"B9",X"05",X"CA",X"05",X"DB",X"05",X"E5",X"05",X"F7",X"05",X"0C",X"06",X"20",X"06",X"33",X"06",
		X"46",X"06",X"59",X"06",X"6C",X"06",X"7F",X"06",X"92",X"06",X"A5",X"06",X"B8",X"06",X"CB",X"06",
		X"96",X"4A",X"47",X"41",X"4D",X"45",X"40",X"40",X"4F",X"56",X"45",X"52",X"3F",X"F1",X"4A",X"50",
		X"55",X"53",X"48",X"40",X"53",X"54",X"41",X"52",X"54",X"40",X"42",X"55",X"54",X"54",X"4F",X"4E",
		X"3F",X"94",X"4A",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"4F",X"4E",X"45",X"3F",X"94",X"4A",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"54",X"57",X"4F",X"3F",X"80",X"4A",X"48",X"49",X"47",
		X"48",X"40",X"53",X"43",X"4F",X"52",X"45",X"3F",X"9F",X"4B",X"40",X"43",X"52",X"45",X"44",X"49",
		X"54",X"40",X"40",X"40",X"40",X"40",X"3F",X"51",X"4B",X"48",X"4F",X"57",X"40",X"46",X"41",X"52",
		X"40",X"43",X"41",X"4E",X"40",X"59",X"4F",X"55",X"40",X"49",X"4E",X"56",X"41",X"44",X"45",X"3F",
		X"5E",X"4B",X"46",X"55",X"45",X"4C",X"3F",X"CC",X"4A",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",
		X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",X"53",X"3F",X"6E",X"4B",X"59",X"4F",X"55",X"40",X"43",
		X"4F",X"4D",X"50",X"4C",X"45",X"54",X"45",X"44",X"40",X"59",X"4F",X"55",X"52",X"40",X"44",X"55",
		X"54",X"49",X"45",X"53",X"3F",X"70",X"4B",X"47",X"4F",X"4F",X"44",X"40",X"4C",X"55",X"43",X"4B",
		X"40",X"4E",X"45",X"58",X"54",X"40",X"54",X"49",X"4D",X"45",X"40",X"41",X"47",X"41",X"49",X"4E",
		X"3F",X"26",X"4A",X"50",X"4C",X"41",X"59",X"3F",X"A9",X"4A",X"5B",X"40",X"53",X"43",X"52",X"41",
		X"4D",X"42",X"4C",X"45",X"40",X"5B",X"3F",X"C7",X"4A",X"5B",X"40",X"53",X"43",X"4F",X"52",X"45",
		X"40",X"54",X"41",X"42",X"4C",X"45",X"40",X"5B",X"3F",X"D5",X"4A",X"31",X"40",X"43",X"4F",X"49",
		X"4E",X"40",X"40",X"32",X"40",X"50",X"4C",X"41",X"59",X"3F",X"78",X"4B",X"42",X"4F",X"4E",X"55",
		X"53",X"40",X"4A",X"45",X"54",X"40",X"40",X"46",X"4F",X"52",X"3F",X"58",X"49",X"30",X"30",X"30",
		X"40",X"50",X"54",X"53",X"3F",X"D4",X"4A",X"4F",X"4E",X"45",X"40",X"50",X"4C",X"41",X"59",X"45",
		X"52",X"40",X"4F",X"4E",X"4C",X"59",X"3F",X"F4",X"4A",X"4F",X"4E",X"45",X"40",X"4F",X"52",X"40",
		X"54",X"57",X"4F",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"3F",X"04",X"4B",X"5B",X"40",
		X"53",X"43",X"4F",X"52",X"45",X"40",X"52",X"41",X"4E",X"4B",X"49",X"4E",X"47",X"40",X"5B",X"3F",
		X"E7",X"4A",X"31",X"53",X"54",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",
		X"54",X"53",X"3F",X"E9",X"4A",X"32",X"4E",X"44",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"50",X"54",X"53",X"3F",X"EB",X"4A",X"33",X"52",X"44",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"ED",X"4A",X"34",X"54",X"48",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"EF",X"4A",X"35",X"54",
		X"48",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"F1",
		X"4A",X"36",X"54",X"48",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",
		X"53",X"3F",X"F3",X"4A",X"37",X"54",X"48",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"50",X"54",X"53",X"3F",X"F5",X"4A",X"38",X"54",X"48",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"F7",X"4A",X"39",X"54",X"48",X"40",X"40",X"40",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"F9",X"4A",X"31",X"30",X"54",
		X"48",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"50",X"54",X"53",X"3F",X"A7",X"CA",
		X"AC",X"0C",X"3D",X"CA",X"DE",X"0A",X"3D",X"CA",X"CA",X"0C",X"C3",X"87",X"0C",X"60",X"D1",X"60",
		X"D1",X"00",X"00",X"60",X"D1",X"60",X"D1",X"00",X"00",X"60",X"D1",X"60",X"D1",X"00",X"00",X"60",
		X"D1",X"60",X"D1",X"00",X"00",X"70",X"D1",X"70",X"D1",X"00",X"01",X"60",X"D1",X"60",X"D1",X"00",
		X"01",X"60",X"D1",X"60",X"D1",X"00",X"00",X"78",X"D1",X"78",X"D1",X"00",X"01",X"60",X"D1",X"60",
		X"D1",X"00",X"01",X"48",X"D1",X"48",X"D1",X"00",X"00",X"58",X"D1",X"58",X"D1",X"00",X"01",X"48",
		X"D1",X"48",X"D1",X"00",X"00",X"58",X"D1",X"58",X"D1",X"00",X"01",X"58",X"D1",X"58",X"D1",X"00",
		X"01",X"68",X"D1",X"68",X"D1",X"00",X"01",X"68",X"D1",X"68",X"D1",X"00",X"02",X"78",X"D1",X"78",
		X"D1",X"00",X"01",X"78",X"D1",X"78",X"D1",X"00",X"01",X"88",X"D1",X"88",X"D1",X"00",X"01",X"88",
		X"D1",X"88",X"D1",X"00",X"02",X"98",X"D1",X"98",X"D1",X"00",X"01",X"98",X"D1",X"98",X"D1",X"00",
		X"01",X"90",X"D1",X"90",X"D1",X"00",X"04",X"90",X"D1",X"90",X"D1",X"00",X"04",X"90",X"D1",X"90",
		X"D1",X"00",X"01",X"90",X"D1",X"90",X"D1",X"00",X"00",X"A0",X"D1",X"A0",X"D1",X"00",X"01",X"80",
		X"D1",X"80",X"D1",X"00",X"00",X"90",X"D1",X"90",X"D1",X"00",X"01",X"70",X"D1",X"70",X"D1",X"00",
		X"00",X"80",X"D1",X"80",X"D1",X"00",X"01",X"60",X"D1",X"60",X"D1",X"00",X"00",X"70",X"D1",X"70",
		X"D1",X"00",X"01",X"50",X"D1",X"50",X"D1",X"00",X"00",X"60",X"D1",X"60",X"D1",X"00",X"01",X"50",
		X"D1",X"50",X"D1",X"00",X"00",X"48",X"D1",X"48",X"D1",X"00",X"00",X"58",X"D1",X"58",X"D1",X"00",
		X"01",X"50",X"D1",X"50",X"D1",X"00",X"00",X"50",X"D1",X"50",X"D1",X"00",X"00",X"60",X"D1",X"60",
		X"D1",X"00",X"01",X"58",X"D1",X"58",X"D1",X"00",X"00",X"68",X"D1",X"68",X"D1",X"00",X"01",X"60",
		X"D1",X"60",X"D1",X"00",X"00",X"70",X"D1",X"70",X"D1",X"00",X"01",X"68",X"D1",X"68",X"D1",X"00",
		X"00",X"78",X"D1",X"78",X"D1",X"00",X"01",X"70",X"D1",X"70",X"D1",X"00",X"00",X"80",X"D1",X"80",
		X"D1",X"00",X"01",X"80",X"D1",X"80",X"D1",X"00",X"00",X"80",X"D1",X"80",X"D1",X"00",X"00",X"80",
		X"D1",X"80",X"D1",X"00",X"04",X"80",X"D1",X"80",X"D1",X"00",X"02",X"80",X"D1",X"80",X"D1",X"00",
		X"04",X"80",X"D1",X"80",X"D1",X"00",X"01",X"80",X"D1",X"80",X"D1",X"00",X"01",X"78",X"D1",X"78",
		X"D1",X"00",X"01",X"70",X"D1",X"70",X"D1",X"00",X"02",X"68",X"D1",X"68",X"D1",X"00",X"04",X"60",
		X"D1",X"60",X"D1",X"00",X"01",X"60",X"D1",X"60",X"D1",X"00",X"01",X"58",X"D1",X"58",X"D1",X"00",
		X"00",X"58",X"D1",X"58",X"D1",X"00",X"00",X"60",X"D1",X"60",X"D1",X"00",X"01",X"48",X"D1",X"48",
		X"D1",X"00",X"00",X"48",X"D1",X"48",X"D1",X"00",X"00",X"50",X"D1",X"50",X"D1",X"00",X"01",X"48",
		X"D1",X"48",X"D1",X"00",X"01",X"58",X"D1",X"58",X"D1",X"00",X"01",X"48",X"D1",X"48",X"D1",X"00",
		X"00",X"50",X"D1",X"50",X"D1",X"00",X"01",X"48",X"D1",X"48",X"D1",X"00",X"00",X"60",X"D1",X"60",
		X"D1",X"00",X"01",X"50",X"D1",X"50",X"D1",X"00",X"02",X"40",X"D1",X"40",X"D1",X"00",X"00",X"60",
		X"D1",X"60",X"D1",X"00",X"01",X"40",X"D1",X"40",X"D1",X"00",X"00",X"60",X"D1",X"60",X"D1",X"00",
		X"01",X"40",X"D1",X"40",X"D1",X"00",X"00",X"50",X"D1",X"50",X"D1",X"00",X"01",X"40",X"D1",X"40",
		X"D1",X"00",X"00",X"50",X"D1",X"50",X"D1",X"00",X"01",X"60",X"D1",X"60",X"D1",X"00",X"00",X"60",
		X"D1",X"60",X"D1",X"00",X"02",X"60",X"D1",X"60",X"D1",X"00",X"00",X"60",X"D1",X"60",X"D1",X"00",
		X"02",X"60",X"D1",X"60",X"D1",X"00",X"00",X"60",X"D1",X"60",X"D1",X"00",X"02",X"70",X"D1",X"70",
		X"D1",X"00",X"01",X"60",X"D1",X"60",X"D1",X"00",X"01",X"60",X"D1",X"60",X"D1",X"00",X"00",X"78",
		X"D1",X"78",X"D1",X"00",X"01",X"60",X"D1",X"60",X"D1",X"00",X"01",X"48",X"D1",X"48",X"D1",X"00",
		X"00",X"58",X"D1",X"58",X"D1",X"00",X"01",X"48",X"D1",X"48",X"D1",X"00",X"00",X"58",X"D1",X"58",
		X"D1",X"00",X"01",X"58",X"D1",X"58",X"D1",X"00",X"01",X"68",X"D1",X"68",X"D1",X"00",X"01",X"68",
		X"D1",X"68",X"D1",X"00",X"02",X"78",X"D1",X"78",X"D1",X"00",X"01",X"78",X"D1",X"78",X"D1",X"00",
		X"01",X"88",X"D1",X"88",X"D1",X"00",X"01",X"88",X"D1",X"88",X"D1",X"00",X"02",X"98",X"D1",X"98",
		X"D1",X"00",X"01",X"98",X"D1",X"98",X"D1",X"00",X"01",X"90",X"D1",X"90",X"D1",X"00",X"04",X"90",
		X"D1",X"90",X"D1",X"00",X"04",X"90",X"D1",X"90",X"D1",X"00",X"01",X"90",X"D1",X"90",X"D1",X"00",
		X"00",X"A0",X"D1",X"A0",X"D1",X"00",X"01",X"80",X"D1",X"80",X"D1",X"00",X"00",X"90",X"D1",X"90",
		X"D1",X"00",X"01",X"70",X"D1",X"70",X"D1",X"00",X"00",X"80",X"D1",X"80",X"D1",X"00",X"01",X"60",
		X"D1",X"60",X"D1",X"00",X"00",X"70",X"D1",X"70",X"D1",X"00",X"01",X"50",X"D1",X"50",X"D1",X"00",
		X"00",X"60",X"D1",X"60",X"D1",X"00",X"01",X"50",X"D1",X"50",X"D1",X"00",X"00",X"48",X"D1",X"48",
		X"D1",X"00",X"00",X"58",X"D1",X"58",X"D1",X"00",X"01",X"50",X"D1",X"50",X"D1",X"00",X"00",X"50",
		X"D1",X"50",X"D1",X"00",X"00",X"60",X"D1",X"60",X"D1",X"00",X"01",X"58",X"D1",X"58",X"D1",X"00",
		X"00",X"68",X"D1",X"68",X"D1",X"00",X"01",X"60",X"D1",X"60",X"D1",X"00",X"00",X"70",X"D1",X"70",
		X"D1",X"00",X"01",X"68",X"D1",X"68",X"D1",X"00",X"00",X"78",X"D1",X"78",X"D1",X"00",X"01",X"70",
		X"D1",X"70",X"D1",X"00",X"00",X"80",X"D1",X"80",X"D1",X"00",X"01",X"80",X"D1",X"80",X"D1",X"00",
		X"00",X"80",X"D1",X"80",X"D1",X"00",X"00",X"80",X"D1",X"80",X"D1",X"00",X"04",X"80",X"D1",X"80",
		X"D1",X"00",X"02",X"80",X"D1",X"80",X"D1",X"00",X"04",X"80",X"D1",X"80",X"D1",X"00",X"01",X"80",
		X"D1",X"80",X"D1",X"00",X"01",X"78",X"D1",X"78",X"D1",X"00",X"01",X"70",X"D1",X"70",X"D1",X"00",
		X"02",X"68",X"D1",X"68",X"D1",X"00",X"04",X"60",X"D1",X"60",X"D1",X"00",X"01",X"60",X"D1",X"60",
		X"D1",X"00",X"01",X"58",X"D1",X"58",X"D1",X"00",X"00",X"58",X"D1",X"58",X"D1",X"00",X"00",X"60",
		X"D1",X"60",X"D1",X"00",X"01",X"48",X"D1",X"48",X"D1",X"00",X"00",X"48",X"D1",X"48",X"D1",X"00",
		X"00",X"50",X"D1",X"50",X"D1",X"00",X"01",X"48",X"D1",X"48",X"D1",X"00",X"01",X"58",X"D1",X"58",
		X"D1",X"00",X"01",X"48",X"D1",X"48",X"D1",X"00",X"00",X"50",X"D1",X"50",X"D1",X"00",X"01",X"48",
		X"D1",X"48",X"D1",X"00",X"00",X"60",X"D1",X"60",X"D1",X"00",X"01",X"50",X"D1",X"50",X"D1",X"00",
		X"02",X"40",X"D1",X"40",X"D1",X"00",X"00",X"60",X"D1",X"60",X"D1",X"00",X"01",X"40",X"D1",X"40",
		X"D1",X"00",X"00",X"60",X"D1",X"60",X"D1",X"00",X"01",X"40",X"D1",X"40",X"D1",X"00",X"00",X"50",
		X"D1",X"50",X"D1",X"00",X"01",X"60",X"D1",X"60",X"D1",X"00",X"00",X"60",X"D1",X"60",X"D1",X"00",
		X"00",X"60",X"D1",X"60",X"D1",X"00",X"00",X"60",X"D1",X"60",X"D1",X"00",X"00",X"FF",X"3E",X"05",
		X"CD",X"19",X"04",X"3A",X"02",X"40",X"FE",X"63",X"38",X"02",X"3E",X"63",X"CD",X"02",X"0B",X"47",
		X"E6",X"F0",X"28",X"07",X"0F",X"0F",X"0F",X"0F",X"32",X"9F",X"4A",X"78",X"E6",X"0F",X"32",X"7F",
		X"4A",X"C9",X"47",X"E6",X"0F",X"C6",X"00",X"27",X"4F",X"78",X"E6",X"F0",X"28",X"0B",X"0F",X"0F",
		X"0F",X"0F",X"47",X"AF",X"C6",X"16",X"27",X"10",X"FB",X"81",X"27",X"C9",X"3A",X"10",X"41",X"0F",
		X"D0",X"3A",X"30",X"42",X"0F",X"D0",X"2A",X"35",X"42",X"7D",X"E6",X"E0",X"6F",X"11",X"05",X"00",
		X"19",X"3E",X"10",X"06",X"19",X"D7",X"11",X"07",X"00",X"19",X"06",X"19",X"D7",X"DD",X"21",X"30",
		X"42",X"DD",X"7E",X"01",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"77",X"7D",X"E6",X"1F",X"47",X"3E",
		X"1D",X"90",X"28",X"10",X"47",X"0E",X"39",X"3A",X"1D",X"41",X"E6",X"1C",X"28",X"02",X"0E",X"3D",
		X"23",X"71",X"10",X"FC",X"DD",X"7E",X"04",X"DD",X"6E",X"05",X"DD",X"66",X"06",X"77",X"7D",X"E6",
		X"1F",X"47",X"3E",X"1D",X"90",X"28",X"10",X"47",X"0E",X"39",X"3A",X"1D",X"41",X"E6",X"1C",X"28",
		X"02",X"0E",X"D0",X"23",X"71",X"10",X"FC",X"DD",X"36",X"00",X"00",X"DD",X"CB",X"08",X"46",X"C8",
		X"DD",X"7E",X"09",X"DD",X"6E",X"0A",X"DD",X"66",X"0B",X"77",X"7D",X"E6",X"1F",X"D6",X"05",X"28",
		X"10",X"47",X"0E",X"39",X"3A",X"1D",X"41",X"E6",X"1C",X"28",X"02",X"0E",X"D0",X"2B",X"71",X"10",
		X"FC",X"DD",X"7E",X"0C",X"DD",X"6E",X"0D",X"DD",X"66",X"0E",X"77",X"7D",X"E6",X"1F",X"D6",X"05",
		X"28",X"10",X"47",X"0E",X"39",X"3A",X"1D",X"41",X"E6",X"1C",X"28",X"02",X"0E",X"3D",X"2B",X"71",
		X"10",X"FC",X"DD",X"36",X"08",X"00",X"C9",X"11",X"04",X"00",X"06",X"08",X"DD",X"21",X"60",X"42",
		X"D9",X"CD",X"EA",X"0B",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"DD",
		X"7E",X"01",X"87",X"87",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"77",X"3C",X"23",X"77",X"3C",X"11",
		X"1F",X"00",X"19",X"77",X"3C",X"23",X"77",X"DD",X"36",X"00",X"00",X"C9",X"3A",X"05",X"41",X"0F",
		X"4F",X"E6",X"78",X"0F",X"0F",X"0F",X"47",X"3E",X"0F",X"90",X"21",X"BE",X"4A",X"11",X"E0",X"FF",
		X"04",X"05",X"28",X"05",X"36",X"CB",X"19",X"10",X"FB",X"47",X"79",X"E6",X"07",X"D9",X"21",X"41",
		X"0C",X"5F",X"16",X"00",X"19",X"7E",X"D9",X"77",X"04",X"05",X"C8",X"19",X"36",X"3C",X"10",X"FB",
		X"C9",X"3C",X"C4",X"C5",X"C6",X"C7",X"C8",X"C9",X"CA",X"CD",X"0C",X"0C",X"3A",X"01",X"41",X"21",
		X"64",X"4B",X"11",X"E0",X"FF",X"47",X"3E",X"18",X"90",X"04",X"05",X"28",X"05",X"36",X"0C",X"19",
		X"10",X"FB",X"47",X"A7",X"28",X"05",X"36",X"10",X"19",X"10",X"FB",X"3A",X"02",X"41",X"21",X"63",
		X"4B",X"47",X"3E",X"18",X"90",X"04",X"05",X"28",X"05",X"36",X"0D",X"19",X"10",X"FB",X"47",X"A7",
		X"C8",X"36",X"10",X"19",X"10",X"FB",X"C9",X"21",X"BF",X"4B",X"11",X"E0",X"FF",X"06",X"0C",X"36",
		X"10",X"19",X"10",X"FB",X"21",X"BF",X"4B",X"3A",X"08",X"41",X"A7",X"C8",X"FE",X"07",X"38",X"02",
		X"3E",X"06",X"47",X"36",X"0A",X"19",X"36",X"0B",X"19",X"10",X"F8",X"C9",X"3A",X"00",X"41",X"E6",
		X"0F",X"3C",X"47",X"3E",X"10",X"90",X"21",X"5F",X"48",X"11",X"20",X"00",X"36",X"0E",X"19",X"10",
		X"FB",X"A7",X"C8",X"36",X"10",X"19",X"3D",X"20",X"FA",X"C9",X"DD",X"21",X"63",X"4B",X"11",X"E0",
		X"FF",X"21",X"0B",X"0D",X"06",X"18",X"7E",X"DD",X"77",X"00",X"23",X"DD",X"19",X"10",X"F7",X"21",
		X"64",X"4B",X"11",X"E0",X"FF",X"DD",X"21",X"23",X"0D",X"06",X"18",X"DD",X"7E",X"00",X"77",X"DD",
		X"23",X"19",X"10",X"F7",X"3A",X"1E",X"41",X"3C",X"47",X"21",X"64",X"4B",X"36",X"81",X"19",X"36",
		X"82",X"19",X"36",X"82",X"19",X"36",X"83",X"19",X"10",X"F2",X"C9",X"50",X"51",X"52",X"6D",X"53",
		X"54",X"55",X"6D",X"56",X"57",X"55",X"6D",X"58",X"59",X"5A",X"6D",X"5B",X"59",X"5A",X"6D",X"64",
		X"65",X"51",X"66",X"6E",X"6F",X"6F",X"80",X"6E",X"6F",X"6F",X"80",X"6E",X"6F",X"6F",X"80",X"6E",
		X"6F",X"6F",X"80",X"6E",X"6F",X"6F",X"80",X"6E",X"6F",X"6F",X"80",X"6E",X"6F",X"6F",X"80",X"6E",
		X"6F",X"6F",X"80",X"F5",X"C5",X"D5",X"E5",X"08",X"D9",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",
		X"E5",X"AF",X"32",X"01",X"68",X"21",X"20",X"40",X"11",X"00",X"50",X"01",X"80",X"00",X"ED",X"B0",
		X"3A",X"00",X"70",X"3A",X"15",X"40",X"32",X"16",X"40",X"3A",X"13",X"40",X"32",X"15",X"40",X"2A",
		X"10",X"40",X"22",X"13",X"40",X"21",X"12",X"40",X"3A",X"02",X"81",X"2F",X"77",X"2B",X"3A",X"01",
		X"81",X"2F",X"77",X"2B",X"3A",X"00",X"81",X"2F",X"77",X"21",X"5F",X"42",X"35",X"CD",X"B9",X"0D",
		X"CD",X"50",X"30",X"21",X"A5",X"0D",X"E5",X"3A",X"05",X"40",X"EF",X"7C",X"0E",X"7D",X"0F",X"B7",
		X"11",X"DE",X"12",X"F6",X"12",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"D9",X"08",X"E1",
		X"D1",X"C1",X"3E",X"01",X"32",X"01",X"68",X"F1",X"C9",X"21",X"18",X"40",X"7E",X"A7",X"28",X"03",
		X"35",X"3E",X"01",X"32",X"02",X"68",X"21",X"10",X"40",X"7E",X"2C",X"2C",X"2C",X"B6",X"2C",X"2C",
		X"2F",X"A6",X"2C",X"E6",X"C4",X"28",X"21",X"47",X"E6",X"C0",X"28",X"05",X"3E",X"06",X"32",X"18",
		X"40",X"CD",X"34",X"0E",X"21",X"02",X"40",X"7E",X"FE",X"63",X"38",X"02",X"36",X"63",X"3A",X"06",
		X"40",X"0F",X"38",X"04",X"11",X"01",X"07",X"FF",X"21",X"03",X"40",X"5E",X"16",X"06",X"1A",X"1C",
		X"73",X"23",X"86",X"3D",X"77",X"3A",X"B0",X"40",X"0F",X"D0",X"2A",X"B1",X"40",X"7E",X"E6",X"07",
		X"20",X"1B",X"EB",X"2A",X"B3",X"40",X"7E",X"FE",X"3F",X"28",X"11",X"23",X"22",X"B3",X"40",X"D6",
		X"30",X"2A",X"B5",X"40",X"77",X"01",X"E0",X"FF",X"09",X"22",X"B5",X"40",X"EB",X"35",X"C0",X"AF",
		X"32",X"B0",X"40",X"C9",X"3A",X"02",X"82",X"CB",X"67",X"28",X"03",X"E6",X"0F",X"C0",X"21",X"02",
		X"40",X"78",X"E6",X"84",X"28",X"0E",X"34",X"3A",X"00",X"40",X"A7",X"C8",X"34",X"3D",X"C8",X"34",
		X"3D",X"C8",X"34",X"C9",X"3A",X"00",X"40",X"2D",X"34",X"A7",X"28",X"08",X"3D",X"28",X"0A",X"3D",
		X"28",X"0C",X"18",X"0F",X"7E",X"FE",X"02",X"18",X"0D",X"7E",X"FE",X"01",X"18",X"08",X"7E",X"FE",
		X"03",X"18",X"03",X"7E",X"FE",X"04",X"D8",X"36",X"00",X"2C",X"34",X"C9",X"2A",X"0B",X"40",X"06",
		X"20",X"3E",X"10",X"D7",X"22",X"0B",X"40",X"21",X"08",X"40",X"35",X"C0",X"2D",X"2D",X"36",X"00",
		X"2D",X"36",X"01",X"AF",X"32",X"0A",X"40",X"21",X"BD",X"0E",X"CD",X"AD",X"0E",X"11",X"04",X"06",
		X"FF",X"11",X"00",X"05",X"FF",X"1E",X"02",X"FF",X"AF",X"32",X"14",X"45",X"C9",X"11",X"20",X"40",
		X"06",X"20",X"EB",X"36",X"00",X"2C",X"1A",X"77",X"2C",X"13",X"10",X"F7",X"C9",X"00",X"05",X"00",
		X"07",X"07",X"01",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"06",X"00",X"05",X"00",
		X"00",X"01",X"01",X"06",X"03",X"03",X"04",X"04",X"04",X"04",X"00",X"00",X"00",X"02",X"02",X"02",
		X"00",X"00",X"00",X"04",X"04",X"04",X"04",X"04",X"06",X"06",X"06",X"06",X"06",X"00",X"05",X"02",
		X"02",X"02",X"02",X"02",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"06",X"06",X"00",X"06",X"06",X"06",X"00",X"05",X"06",
		X"06",X"06",X"06",X"06",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"06",X"00",X"05",X"04",
		X"04",X"04",X"04",X"04",X"02",X"02",X"02",X"02",X"02",X"02",X"06",X"06",X"06",X"06",X"06",X"06",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"06",X"06",X"06",X"06",X"06",X"00",X"05",X"01",
		X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"03",X"03",X"04",X"04",X"05",X"05",X"06",X"06",X"07",
		X"07",X"01",X"01",X"02",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"06",X"21",X"A9",X"11",
		X"E5",X"3A",X"41",X"45",X"EF",X"99",X"0F",X"C7",X"0F",X"07",X"10",X"29",X"10",X"3E",X"10",X"DB",
		X"10",X"04",X"11",X"25",X"11",X"40",X"11",X"8C",X"11",X"3E",X"01",X"32",X"04",X"68",X"3D",X"32",
		X"03",X"68",X"AF",X"32",X"19",X"40",X"21",X"20",X"40",X"11",X"21",X"40",X"01",X"7F",X"00",X"36",
		X"00",X"ED",X"B0",X"21",X"02",X"48",X"22",X"0B",X"40",X"21",X"09",X"40",X"36",X"20",X"21",X"41",
		X"45",X"34",X"AF",X"32",X"06",X"40",X"C9",X"2A",X"0B",X"40",X"06",X"1E",X"3E",X"10",X"D7",X"11",
		X"02",X"00",X"19",X"22",X"0B",X"40",X"21",X"09",X"40",X"35",X"C0",X"21",X"FD",X"0E",X"CD",X"AD",
		X"0E",X"AF",X"32",X"06",X"68",X"32",X"07",X"68",X"21",X"41",X"45",X"34",X"2D",X"36",X"00",X"11",
		X"01",X"07",X"FF",X"11",X"06",X"06",X"FF",X"11",X"12",X"06",X"FF",X"11",X"0F",X"06",X"FF",X"11",
		X"0B",X"06",X"FF",X"1E",X"0C",X"FF",X"C9",X"21",X"40",X"45",X"35",X"C0",X"2C",X"34",X"21",X"3D",
		X"0F",X"CD",X"AD",X"0E",X"11",X"86",X"06",X"FF",X"11",X"92",X"06",X"FF",X"11",X"8B",X"06",X"FF",
		X"11",X"8C",X"06",X"FF",X"11",X"00",X"02",X"FF",X"C9",X"21",X"40",X"45",X"35",X"C0",X"21",X"02",
		X"48",X"22",X"0B",X"40",X"21",X"09",X"40",X"36",X"20",X"21",X"41",X"45",X"34",X"C9",X"2A",X"0B",
		X"40",X"06",X"1A",X"3E",X"10",X"D7",X"11",X"06",X"00",X"19",X"22",X"0B",X"40",X"21",X"09",X"40",
		X"35",X"C0",X"21",X"1D",X"0F",X"CD",X"AD",X"0E",X"11",X"0D",X"06",X"FF",X"21",X"81",X"10",X"11",
		X"60",X"40",X"01",X"18",X"00",X"ED",X"B0",X"21",X"99",X"10",X"22",X"44",X"45",X"21",X"4A",X"4A",
		X"22",X"46",X"45",X"21",X"40",X"45",X"36",X"32",X"2C",X"34",X"2C",X"36",X"0B",X"2C",X"36",X"06",
		X"C9",X"50",X"1C",X"00",X"4A",X"50",X"1E",X"00",X"62",X"50",X"1A",X"06",X"7B",X"50",X"10",X"04",
		X"92",X"50",X"26",X"05",X"A9",X"50",X"33",X"01",X"C2",X"0C",X"0C",X"0C",X"10",X"10",X"05",X"00",
		X"10",X"20",X"24",X"23",X"0C",X"0C",X"0C",X"10",X"10",X"08",X"00",X"10",X"20",X"24",X"23",X"0C",
		X"0C",X"0C",X"10",X"01",X"00",X"00",X"10",X"20",X"24",X"23",X"0C",X"0C",X"0C",X"10",X"01",X"05",
		X"00",X"10",X"20",X"24",X"23",X"0C",X"0C",X"0C",X"10",X"08",X"00",X"00",X"10",X"20",X"24",X"23",
		X"0C",X"0C",X"0C",X"10",X"1D",X"29",X"23",X"24",X"15",X"22",X"29",X"21",X"40",X"45",X"35",X"C0",
		X"36",X"05",X"2A",X"44",X"45",X"7E",X"23",X"22",X"44",X"45",X"2A",X"46",X"45",X"77",X"11",X"E0",
		X"FF",X"19",X"22",X"46",X"45",X"21",X"42",X"45",X"35",X"C0",X"36",X"0B",X"21",X"40",X"45",X"36",
		X"14",X"2C",X"34",X"C9",X"21",X"40",X"45",X"35",X"C0",X"36",X"01",X"2C",X"35",X"2A",X"46",X"45",
		X"11",X"63",X"01",X"19",X"22",X"46",X"45",X"21",X"43",X"45",X"35",X"C0",X"21",X"40",X"45",X"36",
		X"96",X"2C",X"34",X"34",X"C9",X"21",X"40",X"45",X"35",X"C0",X"2C",X"34",X"21",X"60",X"40",X"3E",
		X"10",X"06",X"18",X"D7",X"CD",X"F6",X"18",X"CD",X"17",X"19",X"21",X"BD",X"0E",X"C3",X"AD",X"0E",
		X"21",X"41",X"45",X"34",X"CD",X"CF",X"12",X"CD",X"F5",X"13",X"3E",X"01",X"32",X"19",X"40",X"21",
		X"01",X"00",X"22",X"80",X"43",X"22",X"A0",X"43",X"AF",X"32",X"82",X"43",X"32",X"0D",X"40",X"21",
		X"00",X"41",X"06",X"40",X"D7",X"21",X"B5",X"31",X"11",X"18",X"41",X"7E",X"12",X"23",X"13",X"7E",
		X"12",X"23",X"7E",X"32",X"1D",X"41",X"11",X"02",X"07",X"FF",X"3E",X"20",X"32",X"15",X"41",X"21",
		X"05",X"41",X"36",X"FF",X"2C",X"36",X"05",X"11",X"07",X"06",X"FF",X"C9",X"CD",X"4B",X"1B",X"CD",
		X"37",X"25",X"CD",X"38",X"26",X"CD",X"AA",X"2A",X"CD",X"C0",X"2F",X"21",X"80",X"43",X"7E",X"2C",
		X"B6",X"0F",X"D8",X"21",X"41",X"45",X"36",X"00",X"C9",X"3A",X"02",X"40",X"A7",X"C8",X"21",X"05",
		X"40",X"34",X"AF",X"32",X"0A",X"40",X"C9",X"21",X"47",X"12",X"E5",X"3A",X"0A",X"40",X"EF",X"C5",
		X"11",X"F3",X"11",X"39",X"12",X"AF",X"32",X"19",X"40",X"3E",X"01",X"32",X"04",X"68",X"3D",X"32",
		X"03",X"68",X"21",X"DD",X"0E",X"CD",X"AD",X"0E",X"21",X"60",X"40",X"06",X"40",X"AF",X"D7",X"32",
		X"B0",X"40",X"32",X"06",X"40",X"21",X"02",X"48",X"22",X"0B",X"40",X"21",X"09",X"40",X"36",X"10",
		X"2C",X"34",X"C9",X"2A",X"0B",X"40",X"06",X"1D",X"3E",X"10",X"D7",X"11",X"03",X"00",X"19",X"06",
		X"1D",X"D7",X"19",X"22",X"0B",X"40",X"21",X"09",X"40",X"35",X"C0",X"2C",X"34",X"AF",X"32",X"06",
		X"68",X"32",X"07",X"68",X"32",X"0D",X"40",X"11",X"01",X"07",X"FF",X"11",X"01",X"06",X"FF",X"1E",
		X"16",X"FF",X"1C",X"FF",X"3A",X"17",X"40",X"47",X"E6",X"0F",X"32",X"78",X"49",X"78",X"E6",X"F0",
		X"C8",X"0F",X"0F",X"0F",X"0F",X"32",X"98",X"49",X"C9",X"3A",X"02",X"40",X"A7",X"C8",X"3D",X"11",
		X"18",X"06",X"28",X"01",X"1C",X"FF",X"C9",X"3A",X"11",X"40",X"CB",X"7F",X"C2",X"87",X"12",X"CB",
		X"77",X"C8",X"3A",X"02",X"40",X"FE",X"02",X"D8",X"D6",X"02",X"32",X"02",X"40",X"21",X"00",X"01",
		X"22",X"0D",X"40",X"AF",X"32",X"0A",X"40",X"3E",X"03",X"32",X"05",X"40",X"3E",X"01",X"32",X"06",
		X"40",X"11",X"04",X"06",X"FF",X"CD",X"9D",X"12",X"CD",X"0E",X"31",X"11",X"00",X"04",X"FF",X"3A",
		X"0E",X"40",X"0F",X"D0",X"1C",X"FF",X"C9",X"3A",X"02",X"40",X"A7",X"28",X"0A",X"3D",X"32",X"02",
		X"40",X"21",X"00",X"00",X"C3",X"60",X"12",X"3E",X"01",X"32",X"05",X"40",X"C9",X"AF",X"21",X"00",
		X"41",X"47",X"D7",X"21",X"30",X"42",X"06",X"10",X"D7",X"21",X"60",X"40",X"06",X"40",X"D7",X"21",
		X"60",X"42",X"01",X"02",X"B0",X"DF",X"32",X"19",X"40",X"21",X"00",X"41",X"11",X"01",X"41",X"01",
		X"C0",X"00",X"36",X"00",X"ED",X"B0",X"3A",X"07",X"40",X"32",X"48",X"41",X"32",X"88",X"41",X"21",
		X"C0",X"41",X"11",X"28",X"C9",X"06",X"20",X"72",X"2C",X"73",X"2C",X"10",X"FA",X"C9",X"3A",X"0A",
		X"40",X"EF",X"0E",X"13",X"30",X"13",X"48",X"13",X"D2",X"13",X"FF",X"17",X"62",X"18",X"B1",X"18",
		X"3F",X"19",X"03",X"1A",X"7A",X"1A",X"3A",X"0A",X"40",X"EF",X"0E",X"13",X"30",X"13",X"8D",X"13",
		X"D2",X"13",X"FF",X"17",X"62",X"18",X"8E",X"19",X"C4",X"19",X"03",X"1A",X"7A",X"1A",X"AF",X"32",
		X"19",X"40",X"21",X"60",X"40",X"06",X"40",X"D7",X"21",X"0A",X"40",X"34",X"2D",X"36",X"20",X"21",
		X"00",X"48",X"22",X"0B",X"40",X"CD",X"17",X"19",X"3E",X"01",X"32",X"06",X"40",X"C3",X"CF",X"12",
		X"2A",X"0B",X"40",X"06",X"20",X"3E",X"10",X"D7",X"22",X"0B",X"40",X"21",X"09",X"40",X"35",X"C0",
		X"2C",X"34",X"21",X"BD",X"0E",X"C3",X"AD",X"0E",X"AF",X"32",X"5F",X"42",X"32",X"06",X"68",X"32",
		X"07",X"68",X"32",X"0D",X"40",X"21",X"0A",X"40",X"34",X"2D",X"36",X"96",X"3A",X"0E",X"40",X"0F",
		X"38",X"25",X"11",X"00",X"05",X"FF",X"1E",X"02",X"FF",X"14",X"FF",X"1E",X"04",X"FF",X"11",X"03",
		X"07",X"FF",X"1E",X"00",X"FF",X"21",X"40",X"41",X"11",X"00",X"41",X"01",X"40",X"00",X"ED",X"B0",
		X"2A",X"1D",X"41",X"22",X"18",X"41",X"C9",X"11",X"01",X"05",X"FF",X"18",X"D5",X"AF",X"32",X"5F",
		X"42",X"3A",X"0F",X"40",X"0F",X"30",X"08",X"3E",X"01",X"32",X"06",X"68",X"32",X"07",X"68",X"3E",
		X"01",X"32",X"0D",X"40",X"21",X"0A",X"40",X"34",X"2D",X"36",X"96",X"11",X"00",X"05",X"FF",X"1C",
		X"FF",X"1C",X"FF",X"11",X"03",X"06",X"FF",X"1C",X"FF",X"11",X"03",X"07",X"FF",X"1E",X"00",X"FF",
		X"21",X"80",X"41",X"11",X"00",X"41",X"01",X"40",X"00",X"ED",X"B0",X"2A",X"1D",X"41",X"22",X"18",
		X"41",X"C9",X"21",X"09",X"40",X"35",X"C0",X"36",X"20",X"2C",X"34",X"11",X"82",X"06",X"FF",X"1E",
		X"07",X"FF",X"CD",X"F6",X"18",X"CD",X"17",X"19",X"CD",X"CF",X"12",X"AF",X"32",X"19",X"40",X"21",
		X"60",X"40",X"06",X"40",X"D7",X"21",X"19",X"48",X"11",X"1C",X"00",X"06",X"1E",X"3E",X"36",X"0E",
		X"39",X"77",X"2C",X"71",X"2C",X"71",X"2C",X"71",X"2C",X"71",X"19",X"10",X"F4",X"C9",X"C8",X"2E",
		X"D0",X"36",X"28",X"63",X"28",X"5E",X"00",X"D0",X"36",X"D0",X"2D",X"28",X"5E",X"30",X"63",X"00",
		X"D8",X"36",X"D8",X"36",X"30",X"5E",X"30",X"5E",X"02",X"D8",X"2F",X"E0",X"36",X"38",X"63",X"38",
		X"5E",X"00",X"E0",X"36",X"D8",X"31",X"38",X"5E",X"40",X"63",X"00",X"D0",X"30",X"C8",X"30",X"48",
		X"62",X"48",X"62",X"00",X"C0",X"30",X"B8",X"31",X"48",X"5D",X"50",X"62",X"00",X"B8",X"36",X"B8",
		X"35",X"50",X"5E",X"5F",X"62",X"00",X"B0",X"34",X"B8",X"2C",X"5F",X"5D",X"5F",X"60",X"00",X"C0",
		X"35",X"B8",X"34",X"50",X"60",X"48",X"60",X"00",X"C0",X"2D",X"C8",X"2C",X"48",X"62",X"50",X"62",
		X"00",X"D0",X"36",X"D0",X"2C",X"50",X"60",X"50",X"62",X"00",X"D8",X"2D",X"D8",X"31",X"5F",X"62",
		X"5F",X"60",X"00",X"D0",X"32",X"C8",X"31",X"5F",X"62",X"5F",X"60",X"00",X"C0",X"32",X"C0",X"2F",
		X"50",X"60",X"48",X"60",X"00",X"C8",X"2F",X"C8",X"33",X"48",X"62",X"48",X"60",X"00",X"C8",X"2C",
		X"D0",X"2C",X"40",X"60",X"38",X"60",X"00",X"D0",X"30",X"D0",X"2D",X"38",X"62",X"40",X"62",X"00",
		X"D0",X"31",X"C8",X"34",X"48",X"62",X"48",X"60",X"00",X"C8",X"30",X"C0",X"30",X"40",X"60",X"38",
		X"61",X"00",X"B8",X"30",X"B0",X"30",X"38",X"62",X"40",X"63",X"00",X"B0",X"2C",X"B0",X"30",X"40",
		X"60",X"38",X"61",X"00",X"B0",X"36",X"B0",X"2C",X"30",X"60",X"30",X"62",X"00",X"B8",X"2C",X"B8",
		X"30",X"38",X"62",X"38",X"60",X"00",X"B8",X"2C",X"C0",X"2C",X"30",X"60",X"30",X"62",X"00",X"C8",
		X"36",X"C0",X"30",X"38",X"62",X"40",X"5C",X"00",X"C0",X"2C",X"C8",X"35",X"38",X"60",X"30",X"61",
		X"00",X"C0",X"30",X"C0",X"2C",X"28",X"5E",X"28",X"60",X"00",X"C0",X"31",X"B8",X"30",X"28",X"62",
		X"30",X"62",X"00",X"B0",X"32",X"B0",X"36",X"38",X"62",X"40",X"62",X"00",X"B0",X"2E",X"B8",X"2D",
		X"48",X"62",X"50",X"62",X"00",X"C0",X"2E",X"C8",X"2D",X"5F",X"62",X"5F",X"3A",X"00",X"D0",X"36",
		X"D0",X"36",X"5F",X"3A",X"5F",X"60",X"01",X"D0",X"36",X"D0",X"36",X"50",X"3A",X"50",X"3A",X"02",
		X"D0",X"36",X"D0",X"36",X"5F",X"62",X"5F",X"3A",X"01",X"D0",X"36",X"D0",X"36",X"5F",X"3A",X"5F",
		X"3A",X"02",X"D0",X"36",X"D0",X"2E",X"5F",X"3A",X"5F",X"3A",X"00",X"D8",X"36",X"D8",X"36",X"5F",
		X"3A",X"5F",X"60",X"04",X"D8",X"36",X"D8",X"36",X"50",X"60",X"48",X"60",X"04",X"D0",X"32",X"D0",
		X"36",X"40",X"60",X"38",X"60",X"00",X"D0",X"36",X"D0",X"36",X"30",X"3A",X"30",X"3A",X"01",X"C8",
		X"31",X"C0",X"32",X"30",X"3A",X"30",X"3A",X"00",X"C0",X"36",X"C0",X"36",X"30",X"3A",X"30",X"3A",
		X"01",X"B8",X"31",X"B0",X"32",X"30",X"3A",X"30",X"60",X"00",X"B0",X"36",X"B0",X"36",X"28",X"3A",
		X"28",X"3A",X"00",X"B0",X"36",X"B0",X"36",X"28",X"3A",X"28",X"3A",X"00",X"B0",X"2E",X"B8",X"2D",
		X"30",X"62",X"30",X"3A",X"00",X"C0",X"36",X"C0",X"2E",X"30",X"3A",X"30",X"3A",X"00",X"C8",X"36",
		X"C8",X"36",X"38",X"62",X"40",X"62",X"04",X"C8",X"36",X"C8",X"36",X"48",X"62",X"48",X"3A",X"01",
		X"C8",X"2E",X"D0",X"36",X"48",X"3A",X"50",X"62",X"00",X"D0",X"36",X"D0",X"36",X"5F",X"62",X"5F",
		X"3A",X"04",X"D0",X"36",X"D0",X"2D",X"5F",X"3A",X"5F",X"60",X"00",X"D8",X"36",X"D8",X"36",X"50",
		X"60",X"48",X"60",X"01",X"D8",X"36",X"D8",X"36",X"40",X"60",X"38",X"60",X"02",X"D0",X"31",X"C8",
		X"32",X"30",X"60",X"28",X"60",X"00",X"C0",X"31",X"B8",X"30",X"28",X"62",X"30",X"62",X"00",X"B0",
		X"32",X"B0",X"36",X"38",X"62",X"40",X"62",X"00",X"B0",X"2E",X"B8",X"2D",X"48",X"62",X"50",X"62",
		X"00",X"C0",X"2E",X"C8",X"2D",X"5F",X"62",X"5F",X"3A",X"00",X"D0",X"36",X"D0",X"36",X"5F",X"3A",
		X"5F",X"60",X"01",X"D0",X"36",X"D0",X"36",X"50",X"3A",X"50",X"3A",X"01",X"D0",X"36",X"D0",X"36",
		X"5F",X"62",X"5F",X"3A",X"02",X"D0",X"36",X"D0",X"36",X"5F",X"3A",X"5F",X"3A",X"02",X"D0",X"36",
		X"D0",X"2E",X"5F",X"3A",X"5F",X"3A",X"00",X"D8",X"36",X"D8",X"36",X"5F",X"3A",X"5F",X"60",X"01",
		X"D8",X"36",X"D8",X"36",X"50",X"60",X"48",X"60",X"01",X"D0",X"32",X"D0",X"36",X"40",X"60",X"38",
		X"60",X"00",X"D0",X"36",X"D0",X"36",X"30",X"3A",X"30",X"3A",X"04",X"C8",X"31",X"C0",X"32",X"30",
		X"3A",X"30",X"3A",X"00",X"C0",X"36",X"C0",X"36",X"30",X"3A",X"30",X"3A",X"01",X"B8",X"31",X"B0",
		X"32",X"30",X"3A",X"30",X"60",X"00",X"B0",X"36",X"B0",X"36",X"28",X"3A",X"28",X"3A",X"00",X"B0",
		X"36",X"B0",X"36",X"28",X"3A",X"28",X"3A",X"00",X"B0",X"2E",X"B8",X"2D",X"30",X"62",X"30",X"3A",
		X"00",X"C0",X"36",X"C0",X"2E",X"30",X"3A",X"30",X"3A",X"00",X"C8",X"36",X"C8",X"36",X"38",X"62",
		X"40",X"62",X"04",X"C8",X"36",X"C8",X"36",X"48",X"62",X"48",X"3A",X"04",X"C8",X"2E",X"D0",X"36",
		X"48",X"3A",X"50",X"62",X"00",X"D0",X"36",X"D0",X"36",X"5F",X"62",X"5F",X"3A",X"01",X"D0",X"36",
		X"D0",X"2D",X"5F",X"3A",X"5F",X"60",X"00",X"D8",X"36",X"D8",X"36",X"50",X"60",X"48",X"60",X"04",
		X"D8",X"36",X"D8",X"36",X"40",X"60",X"38",X"60",X"04",X"D0",X"31",X"C8",X"32",X"30",X"60",X"28",
		X"60",X"00",X"C8",X"2C",X"D0",X"2C",X"28",X"62",X"30",X"62",X"00",X"D8",X"2C",X"E0",X"36",X"38",
		X"62",X"40",X"62",X"00",X"E0",X"36",X"E0",X"36",X"48",X"62",X"50",X"62",X"01",X"E0",X"36",X"D8",
		X"34",X"5F",X"5C",X"50",X"60",X"00",X"E0",X"36",X"E0",X"36",X"48",X"60",X"40",X"60",X"02",X"E0",
		X"36",X"E0",X"36",X"38",X"60",X"30",X"60",X"01",X"E0",X"36",X"E0",X"36",X"28",X"5E",X"30",X"62",
		X"01",X"D8",X"34",X"E0",X"36",X"36",X"5C",X"30",X"60",X"00",X"E0",X"36",X"E0",X"36",X"28",X"5E",
		X"30",X"5C",X"04",X"E0",X"36",X"E0",X"36",X"28",X"5E",X"30",X"62",X"01",X"E0",X"36",X"E0",X"36",
		X"38",X"62",X"40",X"62",X"04",X"D8",X"30",X"D0",X"30",X"48",X"62",X"57",X"5C",X"00",X"C8",X"30",
		X"C0",X"30",X"48",X"60",X"40",X"60",X"00",X"B8",X"30",X"B0",X"34",X"38",X"60",X"30",X"60",X"00",
		X"B8",X"2C",X"C0",X"2C",X"28",X"3A",X"28",X"3A",X"00",X"C8",X"2C",X"D0",X"2C",X"28",X"3A",X"28",
		X"3A",X"00",X"D8",X"2C",X"D8",X"34",X"28",X"3A",X"28",X"3A",X"00",X"E0",X"36",X"E0",X"36",X"28",
		X"3A",X"30",X"5C",X"01",X"E0",X"36",X"E0",X"36",X"28",X"3A",X"28",X"3A",X"02",X"D8",X"30",X"D0",
		X"34",X"28",X"3A",X"28",X"3A",X"00",X"D8",X"2C",X"E0",X"36",X"28",X"3A",X"28",X"3A",X"00",X"E0",
		X"36",X"E0",X"36",X"28",X"3A",X"28",X"3A",X"01",X"E0",X"36",X"E0",X"36",X"28",X"3A",X"28",X"3A",
		X"01",X"E0",X"36",X"E0",X"36",X"28",X"3A",X"28",X"3A",X"01",X"E0",X"36",X"D8",X"34",X"28",X"3A",
		X"28",X"3A",X"00",X"E0",X"36",X"E0",X"36",X"28",X"3A",X"28",X"3A",X"04",X"E0",X"36",X"D8",X"30",
		X"28",X"3A",X"28",X"3A",X"00",X"D0",X"30",X"C8",X"30",X"28",X"3A",X"28",X"60",X"00",X"FF",X"21",
		X"09",X"40",X"35",X"C0",X"36",X"0A",X"2C",X"34",X"3E",X"01",X"32",X"19",X"40",X"21",X"01",X"00",
		X"22",X"80",X"43",X"22",X"A0",X"43",X"AF",X"32",X"82",X"43",X"21",X"08",X"41",X"35",X"11",X"03",
		X"07",X"FF",X"21",X"10",X"41",X"11",X"11",X"41",X"01",X"0D",X"00",X"36",X"00",X"ED",X"B0",X"21",
		X"B5",X"31",X"3A",X"1E",X"41",X"47",X"87",X"80",X"5F",X"16",X"00",X"19",X"7E",X"32",X"18",X"41",
		X"23",X"7E",X"32",X"19",X"41",X"23",X"7E",X"32",X"1D",X"41",X"11",X"02",X"07",X"FF",X"3E",X"08",
		X"32",X"15",X"41",X"3E",X"FF",X"32",X"05",X"41",X"3E",X"05",X"32",X"06",X"41",X"11",X"00",X"07",
		X"FF",X"C9",X"CD",X"4B",X"1B",X"CD",X"37",X"25",X"CD",X"38",X"26",X"CD",X"AA",X"2A",X"CD",X"C0",
		X"2F",X"CD",X"1B",X"1B",X"CD",X"7B",X"31",X"CD",X"26",X"1B",X"21",X"80",X"43",X"7E",X"0F",X"38",
		X"19",X"2C",X"7E",X"0F",X"D8",X"21",X"80",X"43",X"11",X"81",X"43",X"36",X"00",X"01",X"A0",X"01",
		X"ED",X"B0",X"21",X"0A",X"40",X"34",X"2D",X"36",X"64",X"C9",X"3A",X"12",X"41",X"FE",X"FF",X"C0",
		X"21",X"80",X"45",X"36",X"96",X"2C",X"36",X"00",X"21",X"0A",X"40",X"36",X"08",X"2D",X"36",X"64",
		X"C9",X"3A",X"08",X"41",X"A7",X"20",X"28",X"CD",X"F6",X"18",X"CD",X"17",X"19",X"11",X"00",X"06",
		X"FF",X"1E",X"02",X"FF",X"3E",X"01",X"32",X"04",X"68",X"3D",X"32",X"03",X"68",X"21",X"C0",X"45",
		X"36",X"96",X"2C",X"36",X"00",X"3E",X"09",X"32",X"0A",X"40",X"AF",X"32",X"19",X"40",X"C9",X"3A",
		X"0E",X"40",X"0F",X"38",X"09",X"21",X"0A",X"40",X"36",X"03",X"2D",X"36",X"32",X"C9",X"21",X"0A",
		X"40",X"34",X"2D",X"36",X"32",X"C9",X"21",X"03",X"48",X"11",X"05",X"00",X"0E",X"20",X"3E",X"10",
		X"06",X"1B",X"77",X"23",X"10",X"FC",X"19",X"0D",X"20",X"F6",X"21",X"2A",X"40",X"06",X"19",X"AF",
		X"77",X"2C",X"77",X"2C",X"10",X"FA",X"C9",X"21",X"80",X"42",X"11",X"81",X"42",X"01",X"A0",X"02",
		X"36",X"00",X"ED",X"B0",X"21",X"60",X"42",X"11",X"61",X"42",X"01",X"1F",X"00",X"36",X"00",X"ED",
		X"B0",X"21",X"60",X"40",X"11",X"61",X"40",X"01",X"3F",X"00",X"36",X"00",X"ED",X"B0",X"C9",X"21",
		X"09",X"40",X"35",X"C0",X"3A",X"08",X"41",X"A7",X"20",X"10",X"3A",X"0E",X"40",X"0F",X"38",X"19",
		X"3E",X"01",X"32",X"05",X"40",X"AF",X"32",X"41",X"45",X"C9",X"3A",X"88",X"41",X"A7",X"20",X"19",
		X"21",X"0A",X"40",X"36",X"03",X"2D",X"36",X"01",X"C9",X"3A",X"88",X"41",X"A7",X"20",X"0A",X"3E",
		X"01",X"32",X"05",X"40",X"AF",X"32",X"41",X"45",X"C9",X"21",X"00",X"41",X"11",X"40",X"41",X"01",
		X"40",X"00",X"ED",X"B0",X"AF",X"32",X"0A",X"40",X"3E",X"04",X"32",X"05",X"40",X"C9",X"3A",X"08",
		X"41",X"A7",X"20",X"28",X"CD",X"F6",X"18",X"CD",X"17",X"19",X"11",X"00",X"06",X"FF",X"1E",X"03",
		X"FF",X"3E",X"01",X"32",X"04",X"68",X"3D",X"32",X"03",X"68",X"21",X"C0",X"45",X"36",X"96",X"2C",
		X"36",X"00",X"3E",X"09",X"32",X"0A",X"40",X"AF",X"32",X"19",X"40",X"C9",X"21",X"0A",X"40",X"34",
		X"2D",X"36",X"64",X"C9",X"21",X"09",X"40",X"35",X"C0",X"3A",X"08",X"41",X"A7",X"20",X"10",X"3A",
		X"48",X"41",X"A7",X"20",X"0A",X"3E",X"01",X"32",X"05",X"40",X"AF",X"32",X"41",X"45",X"C9",X"3A",
		X"48",X"41",X"A7",X"20",X"09",X"21",X"0A",X"40",X"36",X"03",X"2D",X"36",X"01",X"C9",X"21",X"00",
		X"41",X"11",X"80",X"41",X"01",X"40",X"00",X"ED",X"B0",X"AF",X"32",X"0A",X"40",X"3E",X"03",X"32",
		X"05",X"40",X"C9",X"3A",X"81",X"45",X"EF",X"0D",X"1A",X"35",X"1A",X"50",X"1A",X"CD",X"4B",X"1B",
		X"CD",X"37",X"25",X"CD",X"38",X"26",X"CD",X"C0",X"2F",X"21",X"80",X"45",X"35",X"C0",X"36",X"05",
		X"2C",X"34",X"3E",X"01",X"32",X"04",X"68",X"3E",X"00",X"32",X"03",X"68",X"32",X"19",X"40",X"3E",
		X"08",X"32",X"02",X"82",X"C9",X"21",X"80",X"45",X"35",X"C0",X"2C",X"34",X"CD",X"F6",X"18",X"11",
		X"08",X"06",X"FF",X"1C",X"FF",X"1C",X"FF",X"21",X"5D",X"0F",X"CD",X"AD",X"0E",X"C3",X"17",X"19",
		X"21",X"80",X"45",X"35",X"C0",X"21",X"08",X"41",X"34",X"21",X"00",X"41",X"34",X"11",X"00",X"07",
		X"FF",X"AF",X"32",X"5F",X"42",X"21",X"0A",X"40",X"36",X"03",X"2D",X"36",X"0A",X"CD",X"CF",X"12",
		X"AF",X"32",X"1E",X"41",X"21",X"BD",X"0E",X"C3",X"AD",X"0E",X"3A",X"C1",X"45",X"EF",X"84",X"1A",
		X"98",X"1A",X"B7",X"1A",X"21",X"C0",X"45",X"35",X"C0",X"2C",X"34",X"11",X"80",X"06",X"FF",X"1E",
		X"82",X"FF",X"21",X"3D",X"0F",X"C3",X"AD",X"0E",X"CD",X"C5",X"1A",X"7D",X"FE",X"0A",X"28",X"0B",
		X"87",X"87",X"5F",X"16",X"00",X"21",X"2F",X"40",X"19",X"36",X"00",X"11",X"00",X"02",X"FF",X"21",
		X"C0",X"45",X"36",X"80",X"2C",X"34",X"C9",X"21",X"C0",X"45",X"35",X"C0",X"21",X"0A",X"40",X"36",
		X"07",X"2D",X"36",X"64",X"C9",X"01",X"1E",X"00",X"11",X"03",X"00",X"6A",X"DD",X"21",X"A2",X"40",
		X"3A",X"0D",X"40",X"0F",X"30",X"02",X"DD",X"19",X"FD",X"21",X"00",X"42",X"DD",X"7E",X"02",X"FD",
		X"BE",X"02",X"20",X"0F",X"DD",X"7E",X"01",X"FD",X"BE",X"01",X"20",X"07",X"DD",X"7E",X"00",X"FD",
		X"BE",X"00",X"C8",X"30",X"09",X"FD",X"19",X"2C",X"0D",X"0D",X"0D",X"C8",X"18",X"DE",X"7D",X"21",
		X"1D",X"42",X"11",X"20",X"42",X"ED",X"B8",X"6F",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",X"7E",
		X"01",X"FD",X"77",X"01",X"DD",X"7E",X"02",X"FD",X"77",X"02",X"C9",X"3A",X"5F",X"42",X"E6",X"3F",
		X"C0",X"11",X"0C",X"03",X"FF",X"C9",X"3A",X"07",X"41",X"A7",X"C0",X"21",X"A4",X"40",X"3A",X"0D",
		X"40",X"0F",X"30",X"03",X"21",X"A7",X"40",X"7E",X"A7",X"C8",X"CD",X"B0",X"31",X"21",X"08",X"41",
		X"34",X"11",X"03",X"07",X"FF",X"3E",X"01",X"32",X"07",X"41",X"C9",X"CD",X"24",X"1D",X"CD",X"36",
		X"20",X"CD",X"4F",X"1E",X"CD",X"97",X"21",X"CD",X"BF",X"22",X"CD",X"89",X"23",X"CD",X"C8",X"24",
		X"C3",X"29",X"1E",X"DD",X"7E",X"0E",X"A7",X"28",X"05",X"3D",X"DD",X"77",X"0E",X"C9",X"DD",X"6E",
		X"0C",X"DD",X"66",X"0D",X"7E",X"FE",X"FF",X"28",X"15",X"DD",X"77",X"16",X"23",X"7E",X"DD",X"77",
		X"12",X"23",X"7E",X"DD",X"77",X"0E",X"23",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"C9",X"23",X"7E",
		X"DD",X"77",X"0C",X"23",X"7E",X"DD",X"77",X"0D",X"18",X"C9",X"DD",X"E5",X"E1",X"3E",X"07",X"85",
		X"6F",X"DD",X"36",X"0A",X"00",X"DD",X"7E",X"05",X"DD",X"BE",X"03",X"28",X"04",X"38",X"1E",X"18",
		X"56",X"DD",X"7E",X"06",X"DD",X"BE",X"04",X"28",X"0E",X"38",X"06",X"36",X"00",X"2C",X"36",X"01",
		X"C9",X"36",X"00",X"2C",X"36",X"FF",X"C9",X"36",X"00",X"2C",X"36",X"00",X"C9",X"DD",X"7E",X"06",
		X"DD",X"BE",X"04",X"28",X"2C",X"38",X"15",X"36",X"FF",X"2C",X"36",X"01",X"DD",X"7E",X"03",X"DD",
		X"96",X"05",X"47",X"DD",X"7E",X"06",X"DD",X"96",X"04",X"4F",X"18",X"55",X"36",X"FF",X"2C",X"36",
		X"FF",X"DD",X"7E",X"03",X"DD",X"96",X"05",X"47",X"DD",X"7E",X"04",X"DD",X"96",X"06",X"4F",X"18",
		X"40",X"36",X"FF",X"2C",X"36",X"00",X"C9",X"DD",X"7E",X"06",X"DD",X"BE",X"04",X"28",X"2C",X"38",
		X"15",X"36",X"01",X"2C",X"36",X"01",X"DD",X"7E",X"05",X"DD",X"96",X"03",X"47",X"DD",X"7E",X"06",
		X"DD",X"96",X"04",X"4F",X"18",X"1B",X"36",X"01",X"2C",X"36",X"FF",X"DD",X"7E",X"05",X"DD",X"96",
		X"03",X"47",X"DD",X"7E",X"04",X"DD",X"96",X"06",X"4F",X"18",X"06",X"36",X"01",X"2C",X"36",X"00",
		X"C9",X"79",X"B8",X"28",X"16",X"38",X"0B",X"DD",X"36",X"09",X"00",X"CD",X"64",X"1C",X"DD",X"77",
		X"0B",X"C9",X"DD",X"36",X"09",X"01",X"78",X"41",X"4F",X"18",X"F0",X"DD",X"36",X"09",X"01",X"DD",
		X"36",X"0B",X"FF",X"C9",X"AF",X"67",X"68",X"57",X"59",X"06",X"08",X"CB",X"FF",X"07",X"29",X"A7",
		X"ED",X"52",X"38",X"03",X"10",X"F5",X"C9",X"19",X"CB",X"87",X"10",X"EF",X"C9",X"DD",X"7E",X"04",
		X"DD",X"BE",X"06",X"28",X"4A",X"DD",X"7E",X"03",X"DD",X"BE",X"05",X"28",X"58",X"DD",X"CB",X"09",
		X"46",X"28",X"1E",X"DD",X"7E",X"07",X"DD",X"86",X"03",X"DD",X"77",X"03",X"DD",X"7E",X"0B",X"DD",
		X"86",X"0A",X"DD",X"77",X"0A",X"D0",X"DD",X"7E",X"08",X"DD",X"86",X"04",X"DD",X"77",X"04",X"A7",
		X"C9",X"DD",X"7E",X"08",X"DD",X"86",X"04",X"DD",X"77",X"04",X"DD",X"7E",X"0B",X"DD",X"86",X"0A",
		X"DD",X"77",X"0A",X"D0",X"DD",X"7E",X"07",X"DD",X"86",X"03",X"DD",X"77",X"03",X"A7",X"C9",X"DD",
		X"7E",X"03",X"DD",X"BE",X"05",X"28",X"0C",X"30",X"05",X"DD",X"34",X"03",X"A7",X"C9",X"DD",X"35",
		X"03",X"A7",X"C9",X"37",X"C9",X"DD",X"7E",X"04",X"DD",X"BE",X"06",X"30",X"05",X"DD",X"34",X"04",
		X"A7",X"C9",X"DD",X"35",X"04",X"A7",X"C9",X"DD",X"6E",X"13",X"DD",X"66",X"14",X"7E",X"FE",X"80",
		X"20",X"0C",X"23",X"7E",X"DD",X"77",X"13",X"23",X"7E",X"DD",X"77",X"14",X"18",X"E9",X"DD",X"86",
		X"03",X"DD",X"77",X"03",X"23",X"7E",X"DD",X"86",X"04",X"DD",X"77",X"04",X"23",X"DD",X"75",X"13",
		X"DD",X"74",X"14",X"C9",X"DD",X"21",X"10",X"41",X"DD",X"7E",X"05",X"A7",X"20",X"12",X"DD",X"7E",
		X"04",X"DD",X"77",X"05",X"DD",X"7E",X"06",X"E6",X"0F",X"CC",X"44",X"1D",X"DD",X"34",X"06",X"C9",
		X"DD",X"35",X"05",X"C9",X"CD",X"4A",X"1D",X"C3",X"D8",X"1D",X"FD",X"2A",X"18",X"41",X"3E",X"01",
		X"32",X"10",X"41",X"32",X"30",X"42",X"DD",X"7E",X"06",X"2F",X"E6",X"F0",X"47",X"6F",X"26",X"12",
		X"29",X"29",X"E5",X"FD",X"7E",X"02",X"E6",X"F8",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"19",X"22",
		X"35",X"42",X"FD",X"7E",X"03",X"32",X"34",X"42",X"E1",X"1E",X"20",X"19",X"FD",X"7E",X"00",X"E6",
		X"F8",X"0F",X"0F",X"0F",X"5F",X"19",X"22",X"32",X"42",X"FD",X"7E",X"01",X"32",X"31",X"42",X"78",
		X"0F",X"0F",X"5F",X"21",X"C0",X"41",X"19",X"FD",X"7E",X"02",X"77",X"2C",X"36",X"28",X"2C",X"FD",
		X"7E",X"00",X"77",X"2C",X"36",X"28",X"AF",X"32",X"38",X"42",X"32",X"11",X"41",X"2A",X"18",X"41",
		X"1E",X"09",X"FD",X"7E",X"04",X"A7",X"20",X"02",X"1E",X"06",X"19",X"22",X"18",X"41",X"FD",X"7E",
		X"04",X"A7",X"28",X"05",X"FD",X"7E",X"08",X"18",X"03",X"FD",X"7E",X"05",X"32",X"1A",X"41",X"2A",
		X"35",X"42",X"2B",X"2B",X"22",X"1B",X"41",X"C9",X"FD",X"7E",X"04",X"A7",X"C8",X"68",X"26",X"12",
		X"29",X"29",X"E5",X"FD",X"7E",X"06",X"E6",X"F8",X"0F",X"0F",X"0F",X"5F",X"19",X"22",X"3D",X"42",
		X"FD",X"7E",X"07",X"32",X"3C",X"42",X"E1",X"1E",X"20",X"19",X"FD",X"7E",X"04",X"E6",X"F8",X"0F",
		X"0F",X"0F",X"5F",X"19",X"22",X"3A",X"42",X"FD",X"7E",X"05",X"32",X"39",X"42",X"78",X"0F",X"0F",
		X"5F",X"21",X"C0",X"41",X"19",X"2C",X"FD",X"7E",X"06",X"77",X"2C",X"2C",X"FD",X"7E",X"04",X"77",
		X"3E",X"01",X"32",X"11",X"41",X"32",X"38",X"42",X"C9",X"DD",X"21",X"00",X"45",X"11",X"03",X"00",
		X"06",X"04",X"CD",X"3A",X"1E",X"DD",X"19",X"10",X"F9",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"DD",
		X"7E",X"02",X"D6",X"03",X"DD",X"77",X"02",X"FE",X"1F",X"D0",X"DD",X"CB",X"00",X"86",X"C9",X"DD",
		X"21",X"80",X"43",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"EF",X"73",
		X"1E",X"9A",X"1E",X"5C",X"1F",X"8F",X"1F",X"90",X"1F",X"91",X"1F",X"92",X"1F",X"AD",X"1F",X"E6",
		X"1F",X"E7",X"1F",X"DD",X"36",X"03",X"58",X"DD",X"36",X"23",X"58",X"DD",X"36",X"04",X"D0",X"DD",
		X"36",X"24",X"E0",X"21",X"E8",X"1F",X"22",X"8C",X"43",X"21",X"F7",X"1F",X"22",X"AC",X"43",X"DD",
		X"36",X"0E",X"00",X"DD",X"36",X"2E",X"00",X"DD",X"34",X"02",X"21",X"06",X"41",X"35",X"20",X"1B",
		X"3A",X"00",X"41",X"A7",X"28",X"07",X"3D",X"28",X"08",X"36",X"04",X"18",X"06",X"36",X"06",X"18",
		X"02",X"36",X"05",X"2D",X"35",X"20",X"04",X"DD",X"34",X"02",X"C9",X"DD",X"21",X"A0",X"43",X"CD",
		X"63",X"1B",X"DD",X"21",X"80",X"43",X"CD",X"63",X"1B",X"CD",X"CF",X"1E",X"C3",X"25",X"1F",X"3A",
		X"06",X"40",X"0F",X"30",X"1B",X"3A",X"0D",X"40",X"0F",X"38",X"33",X"3A",X"12",X"40",X"06",X"00",
		X"CB",X"67",X"28",X"02",X"CB",X"C0",X"CB",X"77",X"28",X"02",X"CB",X"C8",X"78",X"0F",X"30",X"0E",
		X"DD",X"7E",X"03",X"3D",X"FE",X"38",X"D8",X"DD",X"77",X"03",X"DD",X"35",X"23",X"C9",X"0F",X"D0",
		X"DD",X"7E",X"03",X"3C",X"FE",X"D8",X"D0",X"DD",X"77",X"03",X"DD",X"34",X"23",X"C9",X"3A",X"12",
		X"40",X"06",X"00",X"CB",X"47",X"28",X"02",X"CB",X"C8",X"3A",X"10",X"40",X"CB",X"47",X"28",X"02",
		X"CB",X"C0",X"78",X"18",X"C8",X"3A",X"06",X"40",X"0F",X"30",X"1E",X"3A",X"0D",X"40",X"0F",X"38",
		X"26",X"3A",X"10",X"40",X"07",X"07",X"07",X"30",X"0E",X"DD",X"7E",X"04",X"3C",X"FE",X"D0",X"D0",
		X"DD",X"77",X"04",X"DD",X"34",X"24",X"C9",X"07",X"D0",X"DD",X"7E",X"04",X"3D",X"FE",X"80",X"D8",
		X"DD",X"77",X"04",X"DD",X"35",X"24",X"C9",X"3A",X"11",X"40",X"18",X"D8",X"DD",X"21",X"A0",X"43",
		X"CD",X"63",X"1B",X"DD",X"21",X"80",X"43",X"CD",X"63",X"1B",X"DD",X"34",X"03",X"DD",X"34",X"23",
		X"DD",X"7E",X"03",X"FE",X"F0",X"D8",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",
		X"02",X"06",X"DD",X"36",X"20",X"00",X"DD",X"36",X"21",X"01",X"DD",X"36",X"22",X"06",X"C9",X"C9",
		X"C9",X"C9",X"21",X"06",X"20",X"22",X"8C",X"43",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"0F",X"6F",
		X"21",X"1E",X"20",X"22",X"AC",X"43",X"DD",X"36",X"2E",X"00",X"DD",X"34",X"02",X"3A",X"5F",X"42",
		X"E6",X"03",X"CC",X"DC",X"1F",X"DD",X"21",X"A0",X"43",X"CD",X"63",X"1B",X"DD",X"21",X"80",X"43",
		X"CD",X"63",X"1B",X"3A",X"15",X"41",X"A7",X"20",X"06",X"DD",X"34",X"04",X"DD",X"34",X"24",X"DD",
		X"35",X"0F",X"C0",X"DD",X"36",X"01",X"00",X"DD",X"36",X"21",X"00",X"C9",X"3A",X"17",X"41",X"3C",
		X"E6",X"07",X"32",X"17",X"41",X"C9",X"C9",X"C9",X"06",X"28",X"05",X"06",X"2A",X"05",X"06",X"2C",
		X"05",X"06",X"2E",X"05",X"FF",X"E8",X"1F",X"00",X"27",X"05",X"00",X"29",X"05",X"00",X"2B",X"05",
		X"00",X"2D",X"05",X"FF",X"F7",X"1F",X"04",X"3C",X"10",X"04",X"3D",X"10",X"04",X"3C",X"10",X"04",
		X"3D",X"10",X"04",X"3C",X"10",X"04",X"3D",X"10",X"04",X"3E",X"10",X"FF",X"06",X"20",X"04",X"BC",
		X"10",X"04",X"BD",X"10",X"04",X"BC",X"10",X"04",X"BD",X"10",X"04",X"BC",X"10",X"04",X"BD",X"10",
		X"04",X"BE",X"10",X"FF",X"1E",X"20",X"DD",X"21",X"80",X"42",X"11",X"20",X"00",X"06",X"08",X"D9",
		X"CD",X"49",X"20",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",
		X"D0",X"DD",X"7E",X"02",X"EF",X"69",X"20",X"B2",X"20",X"CA",X"20",X"CB",X"20",X"E5",X"20",X"E6",
		X"20",X"E7",X"20",X"2A",X"21",X"47",X"21",X"48",X"21",X"2A",X"1B",X"41",X"DD",X"75",X"18",X"DD",
		X"74",X"19",X"3A",X"16",X"41",X"E6",X"0F",X"C6",X"F8",X"DD",X"77",X"04",X"7D",X"E6",X"1F",X"07",
		X"07",X"07",X"C6",X"08",X"DD",X"77",X"03",X"DD",X"7E",X"17",X"A7",X"28",X"15",X"3D",X"28",X"08",
		X"3D",X"28",X"0A",X"21",X"5B",X"21",X"18",X"0D",X"21",X"4F",X"21",X"18",X"08",X"21",X"55",X"21",
		X"18",X"03",X"21",X"49",X"21",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"DD",
		X"34",X"02",X"CD",X"63",X"1B",X"3A",X"15",X"41",X"A7",X"C0",X"DD",X"34",X"04",X"DD",X"7E",X"04",
		X"C6",X"14",X"FE",X"08",X"D0",X"DD",X"36",X"02",X"03",X"C9",X"C9",X"DD",X"6E",X"18",X"DD",X"66",
		X"19",X"3E",X"10",X"77",X"23",X"77",X"11",X"1F",X"00",X"19",X"77",X"23",X"77",X"AF",X"DD",X"77",
		X"00",X"DD",X"77",X"01",X"C9",X"C9",X"C9",X"DD",X"7E",X"17",X"3D",X"28",X"05",X"3D",X"28",X"09",
		X"18",X"23",X"21",X"76",X"21",X"3E",X"3F",X"18",X"21",X"DD",X"46",X"1A",X"3E",X"4F",X"05",X"28",
		X"05",X"05",X"28",X"07",X"18",X"0A",X"21",X"8B",X"21",X"18",X"0F",X"21",X"91",X"21",X"18",X"0A",
		X"21",X"85",X"21",X"18",X"05",X"21",X"67",X"21",X"3E",X"3F",X"DD",X"75",X"0C",X"DD",X"74",X"0D",
		X"DD",X"36",X"0E",X"00",X"DD",X"77",X"0F",X"DD",X"34",X"02",X"CD",X"63",X"1B",X"DD",X"35",X"0F",
		X"28",X"10",X"3A",X"15",X"41",X"A7",X"C0",X"DD",X"34",X"04",X"DD",X"7E",X"04",X"C6",X"14",X"FE",
		X"08",X"D0",X"DD",X"36",X"02",X"03",X"C9",X"C9",X"C9",X"02",X"1C",X"10",X"FF",X"49",X"21",X"02",
		X"10",X"10",X"FF",X"4F",X"21",X"02",X"33",X"10",X"FF",X"55",X"21",X"00",X"2F",X"06",X"00",X"26",
		X"06",X"00",X"1F",X"06",X"FF",X"5B",X"21",X"02",X"38",X"10",X"02",X"39",X"10",X"02",X"3A",X"10",
		X"02",X"3B",X"10",X"FF",X"67",X"21",X"02",X"38",X"10",X"02",X"39",X"10",X"02",X"3A",X"10",X"02",
		X"3B",X"10",X"FF",X"76",X"21",X"02",X"11",X"50",X"FF",X"85",X"21",X"02",X"12",X"50",X"FF",X"8B",
		X"21",X"02",X"13",X"50",X"FF",X"91",X"21",X"DD",X"21",X"C0",X"43",X"11",X"20",X"00",X"06",X"02",
		X"D9",X"CD",X"AA",X"21",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",
		X"0F",X"D0",X"DD",X"7E",X"02",X"EF",X"CA",X"21",X"F3",X"21",X"07",X"22",X"08",X"22",X"09",X"22",
		X"0A",X"22",X"0B",X"22",X"1F",X"22",X"35",X"22",X"36",X"22",X"3A",X"83",X"43",X"C6",X"04",X"DD",
		X"77",X"03",X"3A",X"84",X"43",X"C6",X"08",X"DD",X"77",X"04",X"21",X"37",X"22",X"DD",X"75",X"0C",
		X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"21",X"5E",X"22",X"DD",X"75",X"13",X"DD",X"74",X"14",
		X"DD",X"34",X"02",X"CD",X"63",X"1B",X"CD",X"F7",X"1C",X"DD",X"7E",X"03",X"FE",X"F0",X"D8",X"AF",
		X"DD",X"77",X"00",X"DD",X"77",X"01",X"C9",X"C9",X"C9",X"C9",X"C9",X"21",X"4F",X"22",X"DD",X"75",
		X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"0F",X"23",X"DD",X"34",X"02",X"CD",
		X"63",X"1B",X"DD",X"35",X"0F",X"20",X"05",X"AF",X"DD",X"77",X"01",X"C9",X"3A",X"15",X"41",X"A7",
		X"C0",X"DD",X"34",X"04",X"C9",X"C9",X"C9",X"06",X"21",X"04",X"06",X"22",X"04",X"06",X"21",X"04",
		X"06",X"22",X"04",X"06",X"23",X"08",X"06",X"24",X"08",X"06",X"25",X"FE",X"FF",X"37",X"22",X"06",
		X"38",X"09",X"06",X"39",X"09",X"06",X"3A",X"09",X"06",X"3B",X"09",X"FF",X"4F",X"22",X"00",X"00",
		X"01",X"00",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",
		X"01",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"01",X"FF",X"00",X"FF",X"00",X"FF",X"01",X"FF",
		X"00",X"FF",X"01",X"FF",X"01",X"FF",X"00",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"00",
		X"01",X"00",X"01",X"FF",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",X"00",
		X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"80",X"B4",X"22",X"3A",
		X"1D",X"41",X"A7",X"28",X"03",X"FE",X"08",X"C0",X"DD",X"21",X"00",X"44",X"11",X"20",X"00",X"06",
		X"04",X"D9",X"CD",X"DB",X"22",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",
		X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"EF",X"FB",X"22",X"14",X"23",X"40",X"23",X"40",X"23",X"40",
		X"23",X"40",X"23",X"41",X"23",X"55",X"23",X"6B",X"23",X"6B",X"23",X"21",X"6C",X"23",X"DD",X"75",
		X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"21",X"84",X"23",X"DD",X"75",X"13",X"DD",X"74",
		X"14",X"DD",X"34",X"02",X"CD",X"63",X"1B",X"CD",X"F7",X"1C",X"3A",X"17",X"41",X"DD",X"77",X"16",
		X"3A",X"15",X"41",X"A7",X"20",X"03",X"DD",X"34",X"04",X"DD",X"7E",X"04",X"FE",X"F0",X"38",X"08",
		X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"C9",X"DD",X"7E",X"03",X"FE",X"28",X"D0",X"18",X"F0",
		X"C9",X"21",X"75",X"23",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"DD",X"36",
		X"0F",X"3F",X"DD",X"34",X"02",X"CD",X"63",X"1B",X"DD",X"35",X"0F",X"20",X"05",X"AF",X"DD",X"77",
		X"01",X"C9",X"3A",X"15",X"41",X"A7",X"C0",X"DD",X"34",X"04",X"C9",X"C9",X"00",X"1D",X"10",X"00",
		X"1E",X"10",X"FF",X"6C",X"23",X"06",X"38",X"05",X"06",X"39",X"05",X"06",X"3A",X"05",X"06",X"3B",
		X"05",X"FF",X"75",X"23",X"FF",X"00",X"80",X"84",X"23",X"3A",X"1D",X"41",X"FE",X"02",X"C0",X"DD",
		X"21",X"00",X"44",X"11",X"20",X"00",X"06",X"04",X"D9",X"CD",X"A2",X"23",X"D9",X"DD",X"19",X"10",
		X"F7",X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"EF",X"C2",X"23",
		X"DB",X"23",X"EF",X"23",X"EF",X"23",X"F0",X"23",X"F0",X"23",X"F1",X"23",X"05",X"24",X"1B",X"24",
		X"1B",X"24",X"21",X"1C",X"24",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"21",
		X"31",X"24",X"DD",X"75",X"13",X"DD",X"74",X"14",X"DD",X"34",X"02",X"CD",X"63",X"1B",X"CD",X"F7",
		X"1C",X"DD",X"7E",X"04",X"FE",X"F0",X"D8",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"C9",X"C9",
		X"C9",X"21",X"22",X"24",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"DD",X"36",
		X"0F",X"2B",X"DD",X"34",X"02",X"CD",X"63",X"1B",X"DD",X"35",X"0F",X"20",X"05",X"AF",X"DD",X"77",
		X"01",X"C9",X"3A",X"15",X"41",X"A7",X"C0",X"DD",X"34",X"04",X"C9",X"C9",X"05",X"1A",X"10",X"FF",
		X"1C",X"24",X"04",X"38",X"0B",X"04",X"39",X"0B",X"04",X"3A",X"0B",X"04",X"3B",X"0B",X"FF",X"22",
		X"24",X"FF",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",
		X"00",X"FE",X"00",X"FE",X"02",X"FE",X"00",X"FE",X"02",X"FE",X"00",X"FE",X"02",X"FE",X"02",X"FE",
		X"02",X"FE",X"02",X"00",X"02",X"00",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"00",X"02",X"02",X"02",X"00",X"02",X"02",X"02",X"00",X"02",X"02",X"02",
		X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"02",X"02",X"00",X"02",X"00",X"02",
		X"00",X"02",X"02",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"00",X"02",X"02",X"02",X"00",X"02",
		X"02",X"02",X"00",X"02",X"00",X"02",X"02",X"02",X"02",X"02",X"02",X"00",X"02",X"00",X"02",X"00",
		X"02",X"FE",X"02",X"FE",X"02",X"FE",X"02",X"FE",X"02",X"FE",X"00",X"FE",X"02",X"FE",X"00",X"FE",
		X"02",X"FE",X"00",X"FE",X"02",X"FE",X"00",X"FE",X"02",X"FE",X"00",X"FE",X"00",X"FE",X"00",X"FE",
		X"00",X"FE",X"00",X"FE",X"00",X"80",X"31",X"24",X"3A",X"1D",X"41",X"FE",X"01",X"C0",X"DD",X"21",
		X"00",X"44",X"11",X"20",X"00",X"06",X"04",X"D9",X"CD",X"E1",X"24",X"D9",X"DD",X"19",X"10",X"F7",
		X"C9",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"D0",X"DD",X"7E",X"02",X"EF",X"01",X"25",X"DB",
		X"23",X"EF",X"23",X"EF",X"23",X"F0",X"23",X"F0",X"23",X"F1",X"23",X"05",X"24",X"1B",X"24",X"1B",
		X"24",X"21",X"1D",X"25",X"DD",X"75",X"0C",X"DD",X"74",X"0D",X"DD",X"36",X"0E",X"00",X"21",X"32",
		X"25",X"DD",X"75",X"13",X"DD",X"74",X"14",X"DD",X"34",X"02",X"C3",X"DB",X"23",X"00",X"35",X"05",
		X"00",X"36",X"05",X"00",X"37",X"05",X"00",X"30",X"05",X"00",X"37",X"05",X"00",X"36",X"05",X"FF",
		X"1D",X"25",X"00",X"04",X"80",X"32",X"25",X"CD",X"46",X"25",X"CD",X"5B",X"25",X"CD",X"8C",X"25",
		X"CD",X"96",X"25",X"C3",X"E5",X"25",X"21",X"2A",X"40",X"06",X"19",X"3A",X"16",X"41",X"ED",X"44",
		X"4F",X"3A",X"17",X"41",X"71",X"2C",X"77",X"2C",X"10",X"FA",X"C9",X"21",X"60",X"42",X"DD",X"21",
		X"80",X"42",X"11",X"20",X"00",X"06",X"08",X"CD",X"6F",X"25",X"DD",X"19",X"10",X"F9",X"C9",X"DD",
		X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"36",X"00",X"D0",X"36",X"01",X"2C",X"DD",X"7E",X"12",X"77",
		X"2C",X"DD",X"7E",X"18",X"77",X"2C",X"DD",X"7E",X"19",X"77",X"2C",X"C9",X"DD",X"21",X"80",X"43",
		X"FD",X"21",X"60",X"40",X"18",X"12",X"DD",X"21",X"00",X"44",X"FD",X"21",X"70",X"40",X"18",X"08",
		X"DD",X"21",X"80",X"44",X"FD",X"21",X"70",X"40",X"01",X"08",X"04",X"DD",X"7E",X"00",X"DD",X"B6",
		X"01",X"0F",X"30",X"27",X"DD",X"7E",X"16",X"FD",X"77",X"02",X"DD",X"7E",X"03",X"91",X"FD",X"77",
		X"03",X"DD",X"7E",X"04",X"2F",X"91",X"FD",X"77",X"00",X"DD",X"7E",X"12",X"FD",X"77",X"01",X"11",
		X"20",X"00",X"DD",X"19",X"1E",X"04",X"FD",X"19",X"10",X"D1",X"C9",X"FD",X"36",X"00",X"F8",X"FD",
		X"36",X"03",X"F8",X"18",X"EA",X"DD",X"21",X"80",X"40",X"FD",X"21",X"00",X"45",X"06",X"07",X"CD",
		X"FD",X"25",X"11",X"04",X"00",X"DD",X"19",X"1D",X"FD",X"19",X"10",X"F3",X"C9",X"FD",X"CB",X"00",
		X"46",X"28",X"23",X"FD",X"7E",X"02",X"2F",X"DD",X"77",X"01",X"FD",X"7E",X"01",X"C6",X"05",X"DD",
		X"77",X"03",X"3A",X"0F",X"40",X"0F",X"30",X"06",X"3A",X"0D",X"40",X"0F",X"38",X"11",X"DD",X"7E",
		X"03",X"2F",X"DD",X"77",X"03",X"C9",X"DD",X"36",X"01",X"00",X"DD",X"36",X"03",X"00",X"C9",X"DD",
		X"7E",X"03",X"D6",X"0D",X"DD",X"77",X"03",X"C9",X"CD",X"60",X"26",X"CD",X"C4",X"26",X"CD",X"E0",
		X"26",X"CD",X"F6",X"26",X"CD",X"15",X"27",X"CD",X"97",X"29",X"CD",X"65",X"2A",X"CD",X"F7",X"29",
		X"CD",X"8B",X"28",X"CD",X"F2",X"28",X"CD",X"2C",X"29",X"CD",X"68",X"27",X"CD",X"CC",X"27",X"C9",
		X"3A",X"80",X"43",X"0F",X"D0",X"3A",X"1D",X"41",X"FE",X"02",X"C0",X"DD",X"21",X"00",X"44",X"11",
		X"20",X"00",X"06",X"04",X"CD",X"7C",X"26",X"DD",X"19",X"10",X"F9",X"C9",X"DD",X"CB",X"00",X"46",
		X"C8",X"21",X"83",X"43",X"7E",X"DD",X"96",X"03",X"C6",X"06",X"FE",X"0D",X"D0",X"2C",X"7E",X"C6",
		X"04",X"DD",X"96",X"04",X"C6",X"0D",X"FE",X"19",X"D0",X"DD",X"CB",X"00",X"86",X"DD",X"CB",X"01",
		X"C6",X"DD",X"36",X"02",X"06",X"2D",X"2D",X"36",X"06",X"2D",X"36",X"01",X"2D",X"36",X"00",X"21",
		X"A0",X"43",X"36",X"00",X"2C",X"36",X"01",X"DD",X"36",X"17",X"00",X"3E",X"FF",X"32",X"15",X"41",
		X"CD",X"EE",X"30",X"C9",X"3A",X"80",X"43",X"0F",X"D0",X"3A",X"1D",X"41",X"FE",X"01",X"C0",X"DD",
		X"21",X"00",X"44",X"11",X"20",X"00",X"06",X"04",X"CD",X"7C",X"26",X"DD",X"19",X"10",X"F9",X"C9",
		X"3A",X"80",X"43",X"0F",X"D0",X"DD",X"21",X"80",X"42",X"11",X"20",X"00",X"06",X"08",X"CD",X"7C",
		X"26",X"DD",X"19",X"10",X"F9",X"C9",X"3A",X"80",X"43",X"0F",X"D0",X"3A",X"1D",X"41",X"A7",X"28",
		X"03",X"FE",X"08",X"C0",X"DD",X"21",X"00",X"44",X"11",X"20",X"00",X"06",X"04",X"CD",X"7C",X"26",
		X"DD",X"19",X"10",X"F9",X"C9",X"3A",X"80",X"43",X"0F",X"D0",X"3A",X"16",X"41",X"47",X"3A",X"84",
		X"43",X"D6",X"04",X"90",X"E6",X"F8",X"0F",X"0F",X"C6",X"C0",X"6F",X"26",X"41",X"06",X"03",X"3A",
		X"83",X"43",X"C6",X"03",X"5F",X"D6",X"06",X"57",X"7E",X"BB",X"38",X"10",X"2C",X"7E",X"BA",X"30",
		X"0B",X"2C",X"28",X"03",X"10",X"F2",X"C9",X"2E",X"C0",X"10",X"ED",X"C9",X"21",X"80",X"43",X"36",
		X"00",X"2C",X"36",X"01",X"2C",X"36",X"06",X"21",X"A0",X"43",X"36",X"00",X"2C",X"36",X"01",X"3E",
		X"FF",X"32",X"15",X"41",X"CD",X"EE",X"30",X"C9",X"3A",X"1D",X"41",X"FE",X"02",X"C0",X"FD",X"21",
		X"00",X"45",X"06",X"04",X"11",X"20",X"00",X"CD",X"83",X"27",X"FD",X"23",X"FD",X"23",X"FD",X"23",
		X"10",X"F5",X"C9",X"FD",X"CB",X"00",X"46",X"C8",X"DD",X"21",X"00",X"44",X"0E",X"04",X"D9",X"CD",
		X"99",X"27",X"D9",X"DD",X"19",X"0D",X"20",X"F6",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"FD",X"7E",
		X"01",X"DD",X"96",X"03",X"C6",X"03",X"FE",X"07",X"D0",X"FD",X"7E",X"02",X"DD",X"96",X"04",X"C6",
		X"04",X"FE",X"09",X"D0",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"06",
		X"FD",X"36",X"00",X"00",X"11",X"08",X"03",X"FF",X"CD",X"E6",X"30",X"C9",X"FD",X"21",X"00",X"45",
		X"06",X"04",X"11",X"20",X"00",X"CD",X"E1",X"27",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"F5",
		X"C9",X"FD",X"CB",X"00",X"46",X"C8",X"DD",X"21",X"80",X"42",X"0E",X"08",X"D9",X"CD",X"F7",X"27",
		X"D9",X"DD",X"19",X"0D",X"20",X"F6",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"FD",X"7E",X"01",X"DD",
		X"96",X"03",X"C6",X"07",X"FE",X"0F",X"D0",X"FD",X"7E",X"02",X"DD",X"96",X"04",X"C6",X"04",X"FE",
		X"09",X"D0",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"06",X"FD",X"36",
		X"00",X"00",X"DD",X"7E",X"17",X"A7",X"28",X"08",X"3D",X"28",X"0D",X"3D",X"28",X"1D",X"18",X"4E",
		X"11",X"01",X"03",X"FF",X"CD",X"F6",X"30",X"C9",X"21",X"05",X"41",X"7E",X"C6",X"30",X"30",X"02",
		X"3E",X"FF",X"77",X"11",X"03",X"03",X"FF",X"CD",X"C9",X"30",X"C9",X"ED",X"5F",X"E6",X"03",X"A7",
		X"28",X"08",X"3D",X"28",X"05",X"3D",X"28",X"0E",X"18",X"18",X"DD",X"36",X"1A",X"00",X"11",X"05",
		X"03",X"FF",X"CD",X"D1",X"30",X"C9",X"DD",X"36",X"1A",X"01",X"11",X"06",X"03",X"FF",X"CD",X"D1",
		X"30",X"C9",X"DD",X"36",X"1A",X"02",X"11",X"07",X"03",X"FF",X"CD",X"D1",X"30",X"C9",X"11",X"0D",
		X"03",X"FF",X"CD",X"D1",X"30",X"3E",X"FF",X"32",X"12",X"41",X"C9",X"3A",X"1D",X"41",X"A7",X"28",
		X"03",X"FE",X"08",X"C0",X"FD",X"21",X"00",X"45",X"06",X"04",X"11",X"20",X"00",X"CD",X"A9",X"28",
		X"FD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"F5",X"C9",X"FD",X"CB",X"00",X"46",X"C8",X"DD",X"21",
		X"00",X"44",X"0E",X"04",X"D9",X"CD",X"BF",X"28",X"D9",X"DD",X"19",X"0D",X"20",X"F6",X"C9",X"DD",
		X"CB",X"00",X"46",X"C8",X"FD",X"7E",X"01",X"DD",X"96",X"03",X"C6",X"05",X"FE",X"0B",X"D0",X"FD",
		X"7E",X"02",X"DD",X"96",X"04",X"C6",X"03",X"FE",X"07",X"D0",X"DD",X"36",X"00",X"00",X"DD",X"36",
		X"01",X"01",X"DD",X"36",X"02",X"06",X"FD",X"36",X"00",X"00",X"11",X"0A",X"03",X"FF",X"CD",X"F6",
		X"30",X"C9",X"DD",X"21",X"00",X"45",X"11",X"03",X"00",X"06",X"04",X"D9",X"CD",X"05",X"29",X"D9",
		X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"3A",X"16",X"41",X"47",X"DD",X"7E",
		X"02",X"90",X"E6",X"F8",X"0F",X"0F",X"C6",X"C0",X"6F",X"26",X"41",X"7E",X"DD",X"BE",X"01",X"38",
		X"06",X"2C",X"7E",X"DD",X"BE",X"01",X"D8",X"DD",X"36",X"00",X"00",X"C9",X"3A",X"1D",X"41",X"FE",
		X"02",X"C0",X"FD",X"21",X"C0",X"43",X"06",X"02",X"11",X"20",X"00",X"CD",X"43",X"29",X"FD",X"19",
		X"10",X"F9",X"C9",X"FD",X"CB",X"00",X"46",X"C8",X"DD",X"21",X"00",X"44",X"0E",X"04",X"D9",X"CD",
		X"59",X"29",X"D9",X"DD",X"19",X"0D",X"20",X"F6",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"FD",X"7E",
		X"03",X"DD",X"96",X"03",X"C6",X"05",X"FE",X"0B",X"D0",X"FD",X"7E",X"04",X"DD",X"96",X"04",X"C6",
		X"06",X"FE",X"0D",X"D0",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"06",
		X"FD",X"36",X"00",X"00",X"FD",X"36",X"01",X"01",X"FD",X"36",X"02",X"06",X"11",X"08",X"03",X"FF",
		X"CD",X"D9",X"30",X"CD",X"E6",X"30",X"C9",X"FD",X"21",X"C0",X"43",X"06",X"02",X"11",X"20",X"00",
		X"CD",X"A8",X"29",X"FD",X"19",X"10",X"F9",X"C9",X"FD",X"CB",X"00",X"46",X"C8",X"DD",X"21",X"80",
		X"42",X"0E",X"08",X"D9",X"CD",X"BE",X"29",X"D9",X"DD",X"19",X"0D",X"20",X"F6",X"C9",X"DD",X"CB",
		X"00",X"46",X"C8",X"FD",X"7E",X"03",X"DD",X"96",X"03",X"C6",X"07",X"FE",X"0E",X"D0",X"FD",X"7E",
		X"04",X"DD",X"96",X"04",X"C6",X"07",X"FE",X"0E",X"D0",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",
		X"01",X"DD",X"36",X"02",X"06",X"FD",X"36",X"00",X"00",X"FD",X"36",X"01",X"01",X"FD",X"36",X"02",
		X"06",X"CD",X"D9",X"30",X"C3",X"22",X"28",X"3A",X"1D",X"41",X"A7",X"28",X"03",X"FE",X"08",X"C0",
		X"FD",X"21",X"C0",X"43",X"06",X"02",X"11",X"20",X"00",X"CD",X"11",X"2A",X"FD",X"19",X"10",X"F9",
		X"C9",X"FD",X"CB",X"00",X"46",X"C8",X"DD",X"21",X"00",X"44",X"0E",X"04",X"D9",X"CD",X"27",X"2A",
		X"D9",X"DD",X"19",X"0D",X"20",X"F6",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"FD",X"7E",X"03",X"DD",
		X"96",X"03",X"C6",X"06",X"FE",X"0D",X"D0",X"FD",X"7E",X"04",X"DD",X"96",X"04",X"C6",X"04",X"FE",
		X"09",X"D0",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"01",X"DD",X"36",X"02",X"06",X"FD",X"36",
		X"00",X"00",X"FD",X"36",X"01",X"01",X"FD",X"36",X"02",X"06",X"11",X"0A",X"03",X"FF",X"CD",X"D9",
		X"30",X"CD",X"F6",X"30",X"C9",X"DD",X"21",X"C0",X"43",X"06",X"02",X"11",X"20",X"00",X"D9",X"CD",
		X"78",X"2A",X"D9",X"DD",X"19",X"10",X"F7",X"C9",X"DD",X"CB",X"00",X"46",X"C8",X"3A",X"16",X"41",
		X"47",X"DD",X"7E",X"04",X"90",X"E6",X"F8",X"0F",X"0F",X"C6",X"C0",X"6F",X"26",X"41",X"7E",X"DD",
		X"BE",X"03",X"38",X"06",X"2C",X"7E",X"DD",X"BE",X"03",X"D8",X"DD",X"36",X"00",X"00",X"DD",X"36",
		X"01",X"01",X"DD",X"36",X"02",X"06",X"CD",X"D9",X"30",X"C9",X"3A",X"06",X"40",X"0F",X"38",X"19",
		X"3A",X"80",X"43",X"0F",X"30",X"19",X"3A",X"5F",X"42",X"E6",X"67",X"CC",X"0A",X"2B",X"3A",X"5F",
		X"42",X"E6",X"3F",X"CC",X"38",X"2C",X"C3",X"CF",X"2A",X"CD",X"13",X"2C",X"CD",X"E5",X"2A",X"CD",
		X"2D",X"2B",X"CD",X"6A",X"2B",X"CD",X"D6",X"2B",X"CD",X"57",X"2C",X"CD",X"5C",X"2F",X"CD",X"2A",
		X"2F",X"CD",X"8E",X"2F",X"C9",X"3A",X"80",X"43",X"0F",X"D0",X"3A",X"0D",X"40",X"0F",X"38",X"0E",
		X"3A",X"10",X"40",X"CB",X"5F",X"C8",X"3A",X"13",X"40",X"CB",X"5F",X"C0",X"18",X"0C",X"3A",X"11",
		X"40",X"CB",X"5F",X"C8",X"3A",X"14",X"40",X"CB",X"5F",X"C0",X"21",X"00",X"45",X"06",X"04",X"CB",
		X"46",X"20",X"14",X"CB",X"C6",X"2C",X"3A",X"83",X"43",X"C6",X"02",X"77",X"2C",X"3A",X"84",X"43",
		X"D6",X"07",X"77",X"CD",X"FE",X"30",X"C9",X"2C",X"2C",X"2C",X"10",X"E3",X"C9",X"3A",X"1D",X"41",
		X"FE",X"02",X"C0",X"3A",X"5F",X"42",X"E6",X"3F",X"C0",X"DD",X"21",X"00",X"44",X"11",X"20",X"00",
		X"06",X"04",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"30",X"05",X"DD",X"19",X"10",X"F3",X"C9",
		X"DD",X"36",X"00",X"01",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"00",X"DD",X"36",X"03",X"88",
		X"ED",X"5F",X"E6",X"0F",X"C6",X"09",X"DD",X"77",X"04",X"C9",X"3A",X"1D",X"41",X"A7",X"28",X"03",
		X"FE",X"08",X"C0",X"3A",X"5F",X"42",X"E6",X"1F",X"C0",X"ED",X"5F",X"E6",X"01",X"C8",X"DD",X"21",
		X"80",X"42",X"11",X"20",X"00",X"06",X"08",X"DD",X"CB",X"00",X"46",X"20",X"05",X"DD",X"19",X"10",
		X"F6",X"C9",X"DD",X"7E",X"17",X"A7",X"20",X"F5",X"3A",X"A4",X"43",X"DD",X"96",X"04",X"FE",X"70",
		X"30",X"EB",X"FD",X"21",X"00",X"44",X"06",X"04",X"FD",X"7E",X"00",X"FD",X"B6",X"01",X"0F",X"30",
		X"05",X"FD",X"19",X"10",X"F3",X"C9",X"DD",X"36",X"02",X"03",X"DD",X"7E",X"03",X"FD",X"77",X"03",
		X"DD",X"7E",X"04",X"FD",X"77",X"04",X"FD",X"36",X"00",X"01",X"FD",X"36",X"01",X"00",X"FD",X"36",
		X"02",X"00",X"CD",X"08",X"31",X"C9",X"3A",X"1D",X"41",X"FE",X"01",X"C0",X"3A",X"5F",X"42",X"E6",
		X"0F",X"C0",X"DD",X"21",X"00",X"44",X"11",X"20",X"00",X"06",X"04",X"DD",X"7E",X"00",X"DD",X"B6",
		X"01",X"0F",X"30",X"05",X"DD",X"19",X"10",X"F3",X"C9",X"DD",X"36",X"00",X"01",X"DD",X"36",X"01",
		X"00",X"DD",X"36",X"02",X"00",X"ED",X"5F",X"E6",X"7F",X"C6",X"30",X"DD",X"77",X"03",X"DD",X"36",
		X"04",X"08",X"C9",X"3A",X"80",X"43",X"0F",X"D0",X"3A",X"0D",X"40",X"0F",X"38",X"0E",X"3A",X"10",
		X"40",X"CB",X"4F",X"C8",X"3A",X"13",X"40",X"CB",X"4F",X"C0",X"18",X"0C",X"3A",X"11",X"40",X"CB",
		X"57",X"C8",X"3A",X"14",X"40",X"CB",X"57",X"C0",X"21",X"C0",X"43",X"11",X"1F",X"00",X"06",X"02",
		X"7E",X"2C",X"B6",X"0F",X"30",X"04",X"19",X"10",X"F7",X"C9",X"2D",X"36",X"01",X"2C",X"36",X"00",
		X"2C",X"36",X"00",X"CD",X"03",X"31",X"C9",X"3A",X"1A",X"41",X"E6",X"02",X"C8",X"DD",X"21",X"80",
		X"42",X"11",X"20",X"00",X"06",X"08",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",X"30",X"05",X"DD",
		X"19",X"10",X"F3",X"C9",X"DD",X"36",X"00",X"01",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"00",
		X"DD",X"36",X"17",X"01",X"AF",X"32",X"1A",X"41",X"C9",X"C8",X"36",X"CB",X"2E",X"00",X"00",X"D3",
		X"2C",X"DB",X"2E",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"01",X"DB",X"30",X"D3",X"33",X"00",
		X"00",X"D0",X"35",X"CB",X"32",X"00",X"00",X"C3",X"33",X"B8",X"30",X"00",X"00",X"BB",X"2F",X"C3",
		X"2D",X"00",X"00",X"CB",X"2E",X"D3",X"2C",X"00",X"00",X"DB",X"2E",X"E0",X"36",X"00",X"00",X"E0",
		X"36",X"E0",X"36",X"00",X"01",X"E0",X"36",X"E0",X"36",X"00",X"02",X"E0",X"36",X"E0",X"36",X"00",
		X"01",X"DB",X"30",X"D0",X"32",X"00",X"00",X"D3",X"2E",X"DB",X"2C",X"00",X"00",X"DB",X"30",X"D3",
		X"32",X"00",X"00",X"C8",X"34",X"D3",X"2F",X"00",X"00",X"D8",X"36",X"D8",X"36",X"00",X"02",X"D3",
		X"30",X"CB",X"33",X"00",X"00",X"C3",X"30",X"BB",X"33",X"00",X"00",X"B8",X"2F",X"B8",X"30",X"00",
		X"00",X"B8",X"2E",X"C3",X"2D",X"00",X"00",X"CB",X"2C",X"D3",X"2F",X"00",X"00",X"D8",X"36",X"D8",
		X"36",X"00",X"01",X"D8",X"36",X"DB",X"2E",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"04",X"E0",
		X"36",X"E0",X"36",X"00",X"02",X"E0",X"36",X"DB",X"33",X"00",X"00",X"D3",X"30",X"C8",X"30",X"00",
		X"00",X"C0",X"33",X"B8",X"34",X"00",X"00",X"C3",X"2F",X"CB",X"2D",X"00",X"00",X"D3",X"2C",X"DB",
		X"2F",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"02",X"D8",X"32",X"D8",X"35",X"00",X"00",X"DB",
		X"2C",X"E0",X"36",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"04",X"E0",X"36",X"E0",X"36",X"00",
		X"04",X"E0",X"36",X"D8",X"34",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"02",X"E0",X"36",X"E0",
		X"36",X"00",X"01",X"E0",X"36",X"E0",X"36",X"00",X"01",X"D8",X"32",X"D8",X"35",X"00",X"00",X"D0",
		X"30",X"D0",X"2D",X"00",X"00",X"DB",X"2F",X"E0",X"36",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",
		X"04",X"E0",X"36",X"E0",X"36",X"00",X"04",X"E0",X"36",X"E0",X"36",X"00",X"01",X"E0",X"36",X"E0",
		X"36",X"00",X"02",X"E0",X"36",X"E0",X"36",X"00",X"01",X"DB",X"30",X"D3",X"31",X"00",X"00",X"CB",
		X"32",X"C3",X"33",X"00",X"00",X"BB",X"31",X"BB",X"2C",X"00",X"00",X"C3",X"2D",X"CB",X"2E",X"00",
		X"00",X"D0",X"2C",X"D8",X"2E",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"02",X"E0",X"36",X"DB",
		X"33",X"00",X"00",X"D0",X"33",X"CB",X"33",X"00",X"00",X"C8",X"36",X"CB",X"2E",X"00",X"00",X"D3",
		X"2C",X"DB",X"2E",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"04",X"DB",X"30",X"D3",X"33",X"00",
		X"00",X"D0",X"35",X"CB",X"32",X"00",X"00",X"C3",X"33",X"B8",X"30",X"00",X"00",X"BB",X"2F",X"C3",
		X"2D",X"00",X"00",X"CB",X"2E",X"D3",X"2C",X"00",X"00",X"DB",X"2E",X"E0",X"36",X"00",X"00",X"E0",
		X"36",X"E0",X"36",X"00",X"02",X"E0",X"36",X"E0",X"36",X"00",X"01",X"E0",X"36",X"E0",X"36",X"00",
		X"01",X"DB",X"30",X"D0",X"32",X"00",X"00",X"D3",X"2E",X"DB",X"2C",X"00",X"00",X"DB",X"30",X"D3",
		X"32",X"00",X"00",X"C8",X"34",X"D3",X"2F",X"00",X"00",X"D8",X"36",X"D8",X"36",X"00",X"02",X"D3",
		X"30",X"CB",X"33",X"00",X"00",X"C3",X"30",X"BB",X"33",X"00",X"00",X"B8",X"2F",X"B8",X"30",X"00",
		X"00",X"B8",X"2E",X"C3",X"2D",X"00",X"00",X"CB",X"2C",X"D3",X"2F",X"00",X"00",X"D8",X"36",X"D8",
		X"36",X"00",X"00",X"D8",X"36",X"DB",X"2E",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"04",X"E0",
		X"36",X"E0",X"36",X"00",X"02",X"E0",X"36",X"DB",X"33",X"00",X"00",X"D3",X"30",X"C8",X"30",X"00",
		X"00",X"C8",X"36",X"CB",X"2E",X"00",X"00",X"D3",X"2C",X"DB",X"2E",X"00",X"00",X"E0",X"36",X"E0",
		X"36",X"00",X"01",X"DB",X"30",X"D3",X"33",X"00",X"00",X"D0",X"35",X"CB",X"32",X"00",X"00",X"C3",
		X"33",X"B8",X"30",X"00",X"00",X"BB",X"2F",X"C3",X"2D",X"00",X"00",X"CB",X"2E",X"D3",X"2C",X"00",
		X"00",X"DB",X"2E",X"E0",X"36",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"01",X"E0",X"36",X"E0",
		X"36",X"00",X"01",X"E0",X"36",X"E0",X"36",X"00",X"02",X"DB",X"30",X"D0",X"32",X"00",X"00",X"D3",
		X"2E",X"DB",X"2C",X"00",X"00",X"DB",X"30",X"D3",X"32",X"00",X"00",X"C8",X"34",X"D3",X"2F",X"00",
		X"00",X"D8",X"36",X"D8",X"36",X"00",X"02",X"D3",X"30",X"CB",X"33",X"00",X"00",X"C3",X"30",X"BB",
		X"33",X"00",X"00",X"B8",X"2F",X"B8",X"30",X"00",X"00",X"B8",X"2E",X"C3",X"2D",X"00",X"00",X"CB",
		X"2C",X"D3",X"2F",X"00",X"00",X"D8",X"36",X"D8",X"36",X"00",X"00",X"D8",X"36",X"DB",X"2E",X"00",
		X"00",X"E0",X"36",X"E0",X"36",X"00",X"02",X"E0",X"36",X"E0",X"36",X"00",X"04",X"E0",X"36",X"DB",
		X"33",X"00",X"00",X"D3",X"30",X"C8",X"30",X"00",X"00",X"FF",X"3A",X"1A",X"41",X"E6",X"01",X"C8",
		X"DD",X"21",X"80",X"42",X"11",X"20",X"00",X"06",X"08",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"0F",
		X"30",X"05",X"DD",X"19",X"10",X"F3",X"C9",X"DD",X"36",X"00",X"01",X"DD",X"36",X"01",X"00",X"DD",
		X"36",X"02",X"00",X"DD",X"36",X"17",X"00",X"AF",X"32",X"1A",X"41",X"C9",X"3A",X"1A",X"41",X"E6",
		X"04",X"C8",X"DD",X"21",X"80",X"42",X"11",X"20",X"00",X"06",X"08",X"DD",X"7E",X"00",X"DD",X"B6",
		X"01",X"0F",X"30",X"05",X"DD",X"19",X"10",X"F3",X"C9",X"DD",X"36",X"00",X"01",X"DD",X"36",X"01",
		X"00",X"DD",X"36",X"02",X"00",X"DD",X"36",X"17",X"02",X"AF",X"32",X"1A",X"41",X"C9",X"3A",X"1A",
		X"41",X"E6",X"08",X"C8",X"DD",X"21",X"80",X"42",X"11",X"20",X"00",X"06",X"08",X"DD",X"7E",X"00",
		X"DD",X"B6",X"01",X"0F",X"30",X"05",X"DD",X"19",X"10",X"F3",X"C9",X"DD",X"36",X"00",X"01",X"DD",
		X"36",X"01",X"00",X"DD",X"36",X"02",X"00",X"DD",X"36",X"17",X"03",X"AF",X"32",X"1A",X"41",X"C9",
		X"CD",X"C7",X"2F",X"CD",X"02",X"30",X"C9",X"2A",X"18",X"41",X"7E",X"FE",X"FF",X"C0",X"21",X"00",
		X"44",X"11",X"01",X"44",X"01",X"80",X"00",X"36",X"00",X"ED",X"B0",X"21",X"1E",X"41",X"7E",X"FE",
		X"05",X"28",X"01",X"34",X"7E",X"47",X"87",X"80",X"5F",X"16",X"00",X"21",X"B5",X"31",X"19",X"7E",
		X"32",X"18",X"41",X"23",X"7E",X"32",X"19",X"41",X"23",X"7E",X"32",X"1D",X"41",X"11",X"02",X"07",
		X"FF",X"C9",X"3A",X"5F",X"42",X"A7",X"C0",X"21",X"1B",X"40",X"34",X"7E",X"0F",X"D8",X"21",X"17",
		X"41",X"7E",X"3C",X"E6",X"07",X"FE",X"01",X"28",X"03",X"77",X"18",X"02",X"3C",X"77",X"47",X"3A",
		X"11",X"41",X"0F",X"38",X"13",X"78",X"21",X"40",X"30",X"16",X"00",X"87",X"5F",X"19",X"7E",X"32",
		X"04",X"68",X"23",X"7E",X"32",X"03",X"68",X"C9",X"AF",X"32",X"04",X"68",X"32",X"03",X"68",X"C9",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"00",
		X"11",X"41",X"42",X"1A",X"6F",X"26",X"42",X"7E",X"FE",X"FF",X"C8",X"47",X"3A",X"06",X"40",X"A7",
		X"78",X"C4",X"AD",X"30",X"36",X"FF",X"7D",X"FE",X"5E",X"28",X"03",X"3C",X"12",X"C9",X"3E",X"43",
		X"12",X"C9",X"C5",X"D5",X"E5",X"47",X"11",X"40",X"42",X"1A",X"6F",X"26",X"42",X"70",X"7D",X"FE",
		X"5E",X"28",X"04",X"3C",X"12",X"18",X"03",X"3E",X"43",X"12",X"E1",X"D1",X"C1",X"C9",X"3A",X"42",
		X"42",X"F6",X"10",X"32",X"42",X"42",X"32",X"01",X"82",X"AF",X"C3",X"AD",X"30",X"AF",X"CD",X"AD",
		X"30",X"3A",X"42",X"42",X"E6",X"EF",X"32",X"42",X"42",X"32",X"01",X"82",X"C9",X"32",X"00",X"82",
		X"3A",X"42",X"42",X"E6",X"F7",X"32",X"01",X"82",X"00",X"00",X"00",X"00",X"3A",X"42",X"42",X"F6",
		X"08",X"32",X"01",X"82",X"C9",X"3E",X"08",X"18",X"E4",X"3E",X"01",X"CD",X"72",X"30",X"C3",X"31",
		X"31",X"3E",X"01",X"CD",X"72",X"30",X"C3",X"31",X"31",X"3E",X"30",X"CD",X"72",X"30",X"3E",X"02",
		X"CD",X"72",X"30",X"C3",X"31",X"31",X"3E",X"04",X"CD",X"72",X"30",X"C3",X"31",X"31",X"3E",X"05",
		X"CD",X"72",X"30",X"C3",X"31",X"31",X"3E",X"03",X"CD",X"72",X"30",X"C3",X"31",X"31",X"3E",X"06",
		X"C3",X"72",X"30",X"3E",X"20",X"C3",X"72",X"30",X"C9",X"3E",X"0A",X"C3",X"72",X"30",X"3E",X"09",
		X"CD",X"72",X"30",X"3E",X"0A",X"C3",X"72",X"30",X"3E",X"0B",X"CD",X"72",X"30",X"3E",X"0C",X"CD",
		X"72",X"30",X"3E",X"0D",X"C3",X"72",X"30",X"3E",X"0E",X"CD",X"72",X"30",X"3E",X"0F",X"C3",X"72",
		X"30",X"3E",X"13",X"CD",X"72",X"30",X"3E",X"14",X"CD",X"72",X"30",X"3E",X"15",X"C3",X"72",X"30",
		X"3A",X"42",X"42",X"F6",X"40",X"B0",X"32",X"42",X"42",X"32",X"01",X"82",X"C9",X"3A",X"42",X"42",
		X"E6",X"BF",X"32",X"42",X"42",X"32",X"01",X"82",X"AF",X"32",X"1C",X"40",X"C9",X"3E",X"12",X"C3",
		X"72",X"30",X"3E",X"21",X"C3",X"72",X"30",X"3E",X"07",X"C3",X"72",X"30",X"3E",X"22",X"CD",X"72",
		X"30",X"3E",X"23",X"C3",X"72",X"30",X"3E",X"24",X"C3",X"72",X"30",X"3A",X"5F",X"42",X"E6",X"3F",
		X"C0",X"3A",X"05",X"41",X"FE",X"50",X"DC",X"67",X"31",X"3A",X"1D",X"41",X"FE",X"00",X"CC",X"5D",
		X"31",X"FE",X"01",X"CC",X"6C",X"31",X"FE",X"02",X"28",X"0D",X"FE",X"04",X"CC",X"76",X"31",X"FE",
		X"08",X"CC",X"5D",X"31",X"C3",X"5D",X"31",X"3A",X"5F",X"42",X"E6",X"7F",X"CA",X"62",X"31",X"C9",
		X"3E",X"08",X"C3",X"72",X"30",X"C7",X"31",X"00",X"0E",X"14",X"02",X"89",X"2C",X"01",X"ED",X"06",
		X"08",X"B8",X"35",X"04",X"A9",X"39",X"10",X"C0",X"33",X"BC",X"31",X"00",X"00",X"B0",X"32",X"AB",
		X"31",X"00",X"00",X"A0",X"33",X"9B",X"30",X"00",X"00",X"93",X"30",X"8B",X"33",X"00",X"00",X"83",
		X"30",X"7B",X"31",X"00",X"00",X"70",X"32",X"68",X"32",X"00",X"00",X"60",X"34",X"6B",X"2D",X"00",
		X"00",X"73",X"2D",X"7B",X"2E",X"00",X"00",X"80",X"36",X"80",X"36",X"00",X"01",X"83",X"2C",X"83",
		X"30",X"00",X"00",X"80",X"36",X"80",X"36",X"00",X"01",X"80",X"36",X"80",X"36",X"00",X"00",X"80",
		X"36",X"80",X"36",X"00",X"01",X"80",X"36",X"80",X"36",X"00",X"00",X"80",X"36",X"80",X"36",X"00",
		X"01",X"80",X"36",X"80",X"36",X"00",X"01",X"80",X"36",X"80",X"36",X"00",X"01",X"80",X"35",X"80",
		X"35",X"00",X"00",X"80",X"36",X"80",X"36",X"00",X"02",X"83",X"35",X"7B",X"30",X"00",X"00",X"73",
		X"30",X"6B",X"31",X"00",X"00",X"60",X"32",X"60",X"2C",X"00",X"00",X"6B",X"2C",X"73",X"2C",X"00",
		X"00",X"7B",X"2F",X"83",X"2F",X"00",X"00",X"8B",X"2E",X"93",X"2D",X"00",X"00",X"98",X"2E",X"A0",
		X"2E",X"00",X"00",X"AB",X"2D",X"B0",X"2F",X"00",X"00",X"BB",X"2C",X"C3",X"2C",X"00",X"00",X"C8",
		X"36",X"C8",X"2E",X"00",X"00",X"D3",X"2D",X"DB",X"2E",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",
		X"01",X"E0",X"36",X"E0",X"36",X"00",X"01",X"D8",X"32",X"D8",X"35",X"00",X"00",X"DB",X"2C",X"E0",
		X"36",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"02",X"E0",X"36",X"E0",X"36",X"00",X"02",X"E0",
		X"36",X"D8",X"34",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"01",X"E0",X"36",X"E0",X"36",X"00",
		X"01",X"E0",X"36",X"E0",X"36",X"00",X"04",X"D8",X"32",X"D8",X"35",X"00",X"00",X"D0",X"30",X"D0",
		X"2D",X"00",X"00",X"DB",X"2F",X"E0",X"36",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"00",X"E0",
		X"36",X"E0",X"36",X"00",X"01",X"E0",X"36",X"E0",X"36",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",
		X"01",X"E0",X"36",X"E0",X"36",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"01",X"E0",X"36",X"E0",
		X"36",X"00",X"04",X"E0",X"36",X"E0",X"36",X"00",X"02",X"D8",X"30",X"D3",X"30",X"00",X"00",X"D0",
		X"2C",X"D8",X"2E",X"00",X"00",X"E0",X"36",X"E0",X"36",X"00",X"01",X"E0",X"36",X"DB",X"33",X"00",
		X"00",X"D0",X"33",X"CB",X"33",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",X"01",X"C0",X"31",X"C0",
		X"36",X"00",X"00",X"C0",X"36",X"C0",X"36",X"00",X"01",X"B9",X"34",X"C0",X"35",X"00",X"00",X"C0",
		X"36",X"C0",X"36",X"00",X"01",X"B8",X"34",X"B8",X"33",X"00",X"00",X"B8",X"36",X"B8",X"36",X"00",
		X"01",X"B8",X"36",X"B8",X"36",X"00",X"01",X"B0",X"33",X"A8",X"34",X"00",X"00",X"B0",X"36",X"B0",
		X"36",X"00",X"04",X"B0",X"36",X"B0",X"36",X"00",X"02",X"A8",X"33",X"A0",X"32",X"00",X"00",X"A0",
		X"36",X"A0",X"36",X"00",X"01",X"A0",X"36",X"A0",X"36",X"00",X"01",X"98",X"34",X"98",X"30",X"00",
		X"00",X"98",X"2C",X"98",X"33",X"00",X"00",X"98",X"36",X"98",X"36",X"00",X"01",X"98",X"36",X"98",
		X"36",X"00",X"01",X"90",X"34",X"90",X"33",X"00",X"00",X"90",X"36",X"90",X"36",X"00",X"01",X"90",
		X"36",X"90",X"36",X"00",X"01",X"8B",X"32",X"83",X"31",X"00",X"00",X"7B",X"33",X"73",X"34",X"00",
		X"00",X"7B",X"2D",X"83",X"2E",X"00",X"00",X"8B",X"2D",X"93",X"2F",X"00",X"00",X"9B",X"2C",X"A3",
		X"2E",X"00",X"00",X"AB",X"2C",X"B3",X"2D",X"00",X"00",X"B8",X"36",X"B8",X"36",X"00",X"01",X"B8",
		X"36",X"B8",X"36",X"00",X"01",X"B3",X"32",X"AB",X"33",X"00",X"00",X"A0",X"34",X"A0",X"34",X"00",
		X"00",X"A8",X"36",X"A8",X"36",X"00",X"01",X"A3",X"32",X"9B",X"32",X"00",X"00",X"90",X"34",X"98",
		X"35",X"00",X"00",X"98",X"36",X"98",X"36",X"00",X"01",X"93",X"30",X"8B",X"33",X"00",X"00",X"83",
		X"32",X"7B",X"30",X"00",X"00",X"73",X"33",X"6B",X"31",X"00",X"00",X"60",X"34",X"6B",X"2E",X"00",
		X"00",X"70",X"35",X"70",X"2E",X"00",X"00",X"78",X"36",X"78",X"36",X"00",X"01",X"7B",X"2D",X"83",
		X"2D",X"00",X"00",X"88",X"36",X"88",X"36",X"00",X"02",X"8B",X"2F",X"93",X"2D",X"00",X"00",X"9B",
		X"2E",X"A0",X"35",X"00",X"00",X"A0",X"36",X"A0",X"36",X"00",X"01",X"A3",X"2C",X"A3",X"30",X"00",
		X"00",X"9B",X"33",X"90",X"33",X"00",X"00",X"90",X"36",X"90",X"36",X"00",X"01",X"90",X"36",X"90",
		X"36",X"00",X"04",X"88",X"30",X"88",X"2C",X"00",X"00",X"90",X"36",X"90",X"36",X"00",X"01",X"88",
		X"34",X"93",X"2E",X"00",X"00",X"9B",X"2D",X"A3",X"2F",X"00",X"00",X"AB",X"2C",X"B3",X"2E",X"00",
		X"00",X"BB",X"2F",X"C3",X"2C",X"00",X"00",X"C8",X"36",X"CB",X"2E",X"00",X"00",X"D0",X"36",X"D0",
		X"36",X"00",X"01",X"D0",X"35",X"C8",X"34",X"00",X"00",X"D0",X"36",X"D0",X"36",X"00",X"02",X"D0",
		X"36",X"D0",X"36",X"00",X"02",X"CB",X"31",X"C3",X"33",X"00",X"00",X"C0",X"36",X"C0",X"36",X"00",
		X"01",X"C0",X"36",X"BB",X"32",X"00",X"00",X"B0",X"30",X"B0",X"2E",X"00",X"00",X"B8",X"36",X"B3",
		X"33",X"00",X"00",X"AB",X"32",X"AB",X"2C",X"00",X"00",X"B3",X"2C",X"BB",X"2C",X"00",X"00",X"C3",
		X"2C",X"C8",X"36",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",X"01",X"C8",X"36",X"C8",X"35",X"00",
		X"00",X"C8",X"36",X"C0",X"34",X"00",X"00",X"CB",X"2C",X"D3",X"2C",X"00",X"00",X"DB",X"2C",X"DB",
		X"30",X"00",X"00",X"D8",X"36",X"D8",X"36",X"00",X"02",X"DB",X"2D",X"E0",X"36",X"00",X"00",X"E0",
		X"36",X"E0",X"36",X"00",X"04",X"D8",X"34",X"D8",X"30",X"00",X"00",X"D8",X"36",X"D8",X"36",X"00",
		X"01",X"D3",X"30",X"CB",X"32",X"00",X"00",X"C8",X"36",X"C8",X"36",X"00",X"01",X"C8",X"36",X"C8",
		X"36",X"00",X"04",X"CB",X"2C",X"D0",X"35",X"00",X"00",X"CB",X"30",X"C8",X"36",X"00",X"00",X"C0",
		X"33",X"BB",X"33",X"00",X"00",X"B3",X"31",X"AB",X"33",X"00",X"00",X"A0",X"34",X"A8",X"35",X"00",
		X"00",X"A8",X"36",X"A8",X"36",X"00",X"01",X"A8",X"36",X"A8",X"36",X"00",X"01",X"A8",X"36",X"A8",
		X"36",X"00",X"04",X"A8",X"36",X"A8",X"36",X"00",X"02",X"A8",X"35",X"A8",X"2C",X"00",X"00",X"B0",
		X"36",X"B0",X"36",X"00",X"01",X"B0",X"36",X"B0",X"36",X"00",X"01",X"B0",X"36",X"B0",X"36",X"00",
		X"01",X"B0",X"36",X"B0",X"36",X"00",X"00",X"A8",X"34",X"A8",X"31",X"00",X"00",X"A8",X"36",X"A8",
		X"36",X"00",X"02",X"A8",X"36",X"A8",X"36",X"00",X"01",X"A8",X"36",X"A8",X"36",X"00",X"04",X"AB",
		X"2F",X"B3",X"2E",X"00",X"00",X"BB",X"2D",X"C0",X"35",X"00",X"00",X"C0",X"36",X"C0",X"36",X"00",
		X"02",X"BB",X"31",X"B3",X"32",X"00",X"00",X"AB",X"31",X"A0",X"34",X"00",X"00",X"A3",X"31",X"9B",
		X"32",X"00",X"00",X"93",X"33",X"90",X"35",X"00",X"00",X"8B",X"32",X"80",X"34",X"00",X"00",X"8B",
		X"2C",X"93",X"2E",X"00",X"00",X"9B",X"2F",X"A3",X"2C",X"00",X"00",X"AB",X"2D",X"B3",X"2E",X"00",
		X"00",X"BB",X"2D",X"C3",X"2F",X"00",X"00",X"FF",X"60",X"D1",X"60",X"D1",X"47",X"D1",X"47",X"D1",
		X"02",X"60",X"D1",X"60",X"D1",X"47",X"D1",X"47",X"D1",X"02",X"60",X"D1",X"60",X"D1",X"37",X"D1",
		X"37",X"D1",X"00",X"60",X"D1",X"60",X"D1",X"37",X"D1",X"37",X"D1",X"00",X"60",X"D1",X"60",X"D1",
		X"37",X"D1",X"37",X"D1",X"00",X"50",X"D1",X"50",X"D1",X"37",X"D1",X"37",X"D1",X"02",X"50",X"D1",
		X"50",X"D1",X"37",X"D1",X"37",X"D1",X"00",X"60",X"D1",X"60",X"D1",X"37",X"D1",X"37",X"D1",X"00",
		X"60",X"D1",X"60",X"D1",X"37",X"D1",X"37",X"D1",X"00",X"60",X"D1",X"60",X"D1",X"37",X"D1",X"37",
		X"D1",X"00",X"60",X"D1",X"60",X"D1",X"47",X"D1",X"47",X"D1",X"00",X"60",X"D1",X"60",X"D1",X"47",
		X"D1",X"47",X"D1",X"00",X"60",X"D1",X"60",X"D1",X"47",X"D1",X"47",X"D1",X"02",X"60",X"D1",X"60",
		X"D1",X"47",X"D1",X"47",X"D1",X"02",X"60",X"D1",X"60",X"D1",X"47",X"D1",X"47",X"D1",X"02",X"60",
		X"D1",X"60",X"D1",X"2F",X"D1",X"2F",X"D1",X"02",X"60",X"D1",X"60",X"D1",X"2F",X"D1",X"2F",X"D1",
		X"00",X"60",X"D1",X"60",X"D1",X"2F",X"D1",X"2F",X"D1",X"00",X"40",X"D1",X"40",X"D1",X"2F",X"D1",
		X"2F",X"D1",X"00",X"40",X"D1",X"40",X"D1",X"2F",X"D1",X"2F",X"D1",X"00",X"40",X"D1",X"40",X"D1",
		X"2F",X"D1",X"2F",X"D1",X"00",X"40",X"D1",X"40",X"D1",X"2F",X"D1",X"2F",X"D1",X"00",X"40",X"D1",
		X"40",X"D1",X"2F",X"D1",X"2F",X"D1",X"00",X"A0",X"D1",X"A0",X"D1",X"2F",X"D1",X"2F",X"D1",X"00",
		X"A0",X"D1",X"A0",X"D1",X"2F",X"D1",X"2F",X"D1",X"00",X"A0",X"D1",X"A0",X"D1",X"2F",X"D1",X"2F",
		X"D1",X"00",X"A0",X"D1",X"A0",X"D1",X"2F",X"D1",X"2F",X"D1",X"00",X"A0",X"D1",X"A0",X"D1",X"2F",
		X"D1",X"2F",X"D1",X"02",X"A0",X"D1",X"A0",X"D1",X"2F",X"D1",X"2F",X"D1",X"02",X"A0",X"D1",X"A0",
		X"D1",X"37",X"D1",X"37",X"D1",X"02",X"A0",X"D1",X"A0",X"D1",X"8F",X"D1",X"8F",X"D1",X"02",X"A0",
		X"D1",X"A0",X"D1",X"8F",X"D1",X"8F",X"D1",X"02",X"A0",X"D1",X"A0",X"D1",X"8F",X"D1",X"8F",X"D1",
		X"02",X"A0",X"D1",X"A0",X"D1",X"8F",X"D1",X"8F",X"D1",X"00",X"A0",X"D1",X"A0",X"D1",X"8F",X"D1",
		X"8F",X"D1",X"00",X"A0",X"D1",X"A0",X"D1",X"8F",X"D1",X"8F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",
		X"8F",X"D1",X"8F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"8F",X"D1",X"8F",X"D1",X"00",X"D8",X"D1",
		X"D8",X"D1",X"8F",X"D1",X"8F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",X"00",
		X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",X"02",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",
		X"D1",X"02",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",X"02",X"D8",X"D1",X"D8",X"D1",X"C7",
		X"D1",X"C7",X"D1",X"02",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",X"00",X"D8",X"D1",X"D8",
		X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"D8",
		X"D1",X"D8",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"3F",X"D1",X"3F",X"D1",
		X"00",X"D8",X"D1",X"D8",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"3F",X"D1",
		X"3F",X"D1",X"00",X"50",X"D1",X"50",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"50",X"D1",X"50",X"D1",
		X"3F",X"D1",X"3F",X"D1",X"00",X"50",X"D1",X"50",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"50",X"D1",
		X"50",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"50",X"D1",X"50",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",
		X"D8",X"D1",X"D8",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"3F",X"D1",X"3F",
		X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"3F",
		X"D1",X"3F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"D8",X"D1",X"D8",
		X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"D8",
		X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",
		X"00",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",
		X"C7",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",
		X"C7",X"D1",X"C7",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",X"00",X"D8",X"D1",
		X"D8",X"D1",X"4F",X"D1",X"4F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"4F",X"D1",X"4F",X"D1",X"00",
		X"D8",X"D1",X"D8",X"D1",X"4F",X"D1",X"4F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"4F",X"D1",X"4F",
		X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"4F",X"D1",X"4F",X"D1",X"00",X"60",X"D1",X"60",X"D1",X"4F",
		X"D1",X"4F",X"D1",X"00",X"60",X"D1",X"60",X"D1",X"4F",X"D1",X"4F",X"D1",X"00",X"60",X"D1",X"60",
		X"D1",X"4F",X"D1",X"4F",X"D1",X"00",X"60",X"D1",X"60",X"D1",X"37",X"D1",X"37",X"D1",X"00",X"60",
		X"D1",X"60",X"D1",X"37",X"D1",X"37",X"D1",X"00",X"48",X"D1",X"48",X"D1",X"37",X"D1",X"37",X"D1",
		X"00",X"48",X"D1",X"48",X"D1",X"37",X"D1",X"37",X"D1",X"00",X"48",X"D1",X"48",X"D1",X"37",X"D1",
		X"37",X"D1",X"00",X"58",X"D1",X"58",X"D1",X"37",X"D1",X"37",X"D1",X"00",X"58",X"D1",X"58",X"D1",
		X"37",X"D1",X"37",X"D1",X"00",X"58",X"D1",X"58",X"D1",X"47",X"D1",X"47",X"D1",X"00",X"58",X"D1",
		X"58",X"D1",X"47",X"D1",X"47",X"D1",X"00",X"58",X"D1",X"58",X"D1",X"47",X"D1",X"47",X"D1",X"00",
		X"58",X"D1",X"58",X"D1",X"47",X"D1",X"47",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"47",X"D1",X"47",
		X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"47",X"D1",X"47",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"47",
		X"D1",X"47",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"47",X"D1",X"47",X"D1",X"00",X"D8",X"D1",X"D8",
		X"D1",X"47",X"D1",X"47",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",X"00",X"D8",
		X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",
		X"00",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",
		X"C7",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",X"02",X"D8",X"D1",X"D8",X"D1",
		X"C7",X"D1",X"C7",X"D1",X"02",X"D8",X"D1",X"D8",X"D1",X"C7",X"D1",X"C7",X"D1",X"02",X"D8",X"D1",
		X"D8",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",
		X"D8",X"D1",X"D8",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"3F",X"D1",X"3F",
		X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"D8",X"D1",X"D8",X"D1",X"3F",
		X"D1",X"3F",X"D1",X"00",X"50",X"D1",X"50",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"60",X"D1",X"60",
		X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"60",X"D1",X"60",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"60",
		X"D1",X"60",X"D1",X"3F",X"D1",X"3F",X"D1",X"00",X"FF",X"C8",X"D1",X"C8",X"D1",X"00",X"00",X"C8",
		X"D1",X"C8",X"D1",X"00",X"00",X"90",X"D1",X"90",X"D1",X"00",X"00",X"50",X"D1",X"50",X"D1",X"00",
		X"00",X"90",X"D1",X"90",X"D1",X"00",X"00",X"C8",X"D1",X"C8",X"D1",X"00",X"00",X"C8",X"D1",X"C8",
		X"D1",X"00",X"00",X"98",X"D1",X"98",X"D1",X"00",X"00",X"98",X"D1",X"98",X"D1",X"00",X"00",X"98",
		X"D1",X"98",X"D1",X"00",X"00",X"C8",X"D1",X"C8",X"D1",X"00",X"00",X"48",X"D1",X"48",X"D1",X"00",
		X"00",X"48",X"D1",X"48",X"D1",X"00",X"00",X"48",X"D1",X"48",X"D1",X"00",X"00",X"C8",X"D1",X"C8",
		X"D1",X"00",X"00",X"98",X"D1",X"98",X"D1",X"00",X"00",X"98",X"D1",X"98",X"D1",X"00",X"00",X"98",
		X"D1",X"98",X"D1",X"00",X"00",X"C8",X"D1",X"C8",X"D1",X"00",X"00",X"C8",X"D1",X"C8",X"D1",X"00",
		X"00",X"C8",X"D1",X"C8",X"D1",X"00",X"08",X"C8",X"D1",X"C8",X"D1",X"00",X"00",X"C8",X"D1",X"C8",
		X"D1",X"00",X"00",X"C8",X"D1",X"C8",X"D1",X"00",X"00",X"70",X"D1",X"70",X"D1",X"00",X"00",X"70",
		X"D1",X"70",X"D1",X"00",X"00",X"C8",X"D1",X"C8",X"D1",X"00",X"00",X"C8",X"D1",X"C8",X"D1",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
