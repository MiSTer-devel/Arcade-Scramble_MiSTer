library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_SND_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_SND_2 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"88",X"8C",X"8F",X"8C",X"88",X"8C",X"88",X"8C",X"8F",X"8C",X"88",X"AF",X"FF",X"1F",X"0A",X"5F",
		X"09",X"A8",X"80",X"68",X"68",X"A8",X"80",X"68",X"68",X"88",X"83",X"88",X"8C",X"88",X"83",X"88",
		X"83",X"88",X"8C",X"88",X"83",X"88",X"83",X"88",X"8C",X"88",X"83",X"AC",X"FF",X"FF",X"CD",X"C7",
		X"06",X"3E",X"01",X"32",X"73",X"80",X"CD",X"0D",X"05",X"C3",X"8E",X"0F",X"CD",X"C7",X"06",X"CD",
		X"0D",X"05",X"C9",X"CD",X"C7",X"06",X"CD",X"0D",X"05",X"C9",X"DD",X"21",X"50",X"80",X"C3",X"DA",
		X"0D",X"DD",X"21",X"58",X"80",X"C3",X"DA",X"0D",X"DD",X"21",X"60",X"80",X"C3",X"DA",X"0D",X"1F",
		X"0A",X"3F",X"0E",X"5F",X"08",X"85",X"85",X"85",X"8A",X"8A",X"8A",X"8A",X"91",X"91",X"91",X"91",
		X"8F",X"8F",X"D6",X"93",X"8F",X"93",X"B6",X"93",X"8F",X"93",X"B6",X"FF",X"1F",X"0A",X"5F",X"08",
		X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"8E",X"8E",X"8E",X"8E",X"8C",X"8C",X"D3",X"8F",X"8C",
		X"8F",X"B3",X"8F",X"8C",X"8F",X"B3",X"FF",X"1F",X"0A",X"5F",X"08",X"91",X"91",X"91",X"8A",X"8A",
		X"8A",X"8A",X"96",X"96",X"96",X"96",X"94",X"94",X"D6",X"93",X"8F",X"93",X"B6",X"93",X"8F",X"93",
		X"B6",X"FF",X"CD",X"C7",X"06",X"3E",X"02",X"32",X"73",X"80",X"CD",X"0D",X"05",X"C3",X"8E",X"0F",
		X"CD",X"C7",X"06",X"CD",X"0D",X"05",X"C9",X"DD",X"21",X"50",X"80",X"C3",X"DA",X"0D",X"DD",X"21",
		X"58",X"80",X"C3",X"DA",X"0D",X"1F",X"0A",X"3F",X"0A",X"5F",X"09",X"8D",X"8F",X"91",X"8F",X"91",
		X"94",X"91",X"8F",X"8D",X"8F",X"91",X"8D",X"8F",X"8C",X"AD",X"FF",X"1F",X"0A",X"5F",X"09",X"8A",
		X"8C",X"8D",X"8C",X"8D",X"8F",X"8D",X"8C",X"8A",X"8C",X"8D",X"8A",X"8C",X"88",X"AA",X"FF",X"FF",
		X"CD",X"BC",X"07",X"21",X"00",X"03",X"22",X"83",X"80",X"21",X"80",X"80",X"36",X"01",X"21",X"00",
		X"08",X"22",X"81",X"80",X"CD",X"C6",X"04",X"CD",X"0D",X"05",X"06",X"0B",X"CD",X"FE",X"05",X"C9",
		X"2A",X"83",X"80",X"2B",X"22",X"83",X"80",X"7D",X"B4",X"28",X"52",X"3A",X"80",X"80",X"FE",X"00",
		X"28",X"1E",X"FE",X"01",X"28",X"0E",X"FE",X"02",X"28",X"05",X"21",X"00",X"0A",X"18",X"08",X"21",
		X"00",X"06",X"18",X"03",X"21",X"00",X"08",X"22",X"81",X"80",X"CD",X"C6",X"04",X"AF",X"18",X"28",
		X"2A",X"81",X"80",X"11",X"20",X"00",X"ED",X"52",X"22",X"81",X"80",X"7C",X"FE",X"00",X"28",X"06",
		X"CD",X"C6",X"04",X"AF",X"18",X"12",X"CD",X"C6",X"04",X"3A",X"80",X"80",X"3C",X"32",X"80",X"80",
		X"FE",X"04",X"28",X"02",X"AF",X"C9",X"3E",X"01",X"32",X"80",X"80",X"AF",X"C9",X"3E",X"FF",X"C9",
		X"CD",X"BC",X"07",X"3E",X"01",X"32",X"86",X"80",X"3E",X"20",X"32",X"87",X"80",X"3E",X"06",X"32",
		X"88",X"80",X"AF",X"32",X"89",X"80",X"32",X"8A",X"80",X"21",X"00",X"03",X"22",X"8D",X"80",X"21",
		X"00",X"04",X"22",X"8B",X"80",X"CD",X"C6",X"04",X"CD",X"0D",X"05",X"06",X"0B",X"CD",X"FE",X"05",
		X"C9",X"2A",X"8D",X"80",X"2B",X"7C",X"B5",X"28",X"5D",X"22",X"8D",X"80",X"3A",X"89",X"80",X"FE",
		X"00",X"28",X"06",X"FE",X"01",X"28",X"24",X"AF",X"C9",X"21",X"86",X"80",X"35",X"20",X"F8",X"36",
		X"01",X"CD",X"80",X"06",X"B7",X"11",X"08",X"00",X"ED",X"52",X"CD",X"C6",X"04",X"21",X"87",X"80",
		X"35",X"20",X"E4",X"36",X"20",X"21",X"89",X"80",X"34",X"18",X"DC",X"2A",X"8B",X"80",X"11",X"30",
		X"00",X"3A",X"8A",X"80",X"E6",X"01",X"20",X"1B",X"B7",X"ED",X"52",X"22",X"8B",X"80",X"CD",X"C6",
		X"04",X"21",X"88",X"80",X"35",X"20",X"06",X"36",X"06",X"21",X"8A",X"80",X"34",X"21",X"89",X"80",
		X"35",X"18",X"B4",X"19",X"18",X"E5",X"3E",X"FF",X"C9",X"C9",X"3E",X"FF",X"C9",X"CD",X"82",X"07",
		X"3E",X"01",X"32",X"A0",X"80",X"3E",X"20",X"32",X"A1",X"80",X"3E",X"10",X"32",X"A2",X"80",X"AF",
		X"32",X"A5",X"80",X"32",X"A6",X"80",X"21",X"00",X"01",X"22",X"A3",X"80",X"21",X"00",X"05",X"22",
		X"A7",X"80",X"CD",X"C6",X"04",X"CD",X"0D",X"05",X"06",X"0D",X"CD",X"FE",X"05",X"C9",X"2A",X"A3",
		X"80",X"2B",X"7C",X"B5",X"28",X"5D",X"22",X"A3",X"80",X"3A",X"A5",X"80",X"FE",X"00",X"28",X"06",
		X"FE",X"01",X"28",X"24",X"AF",X"C9",X"21",X"A0",X"80",X"35",X"20",X"F8",X"36",X"01",X"CD",X"80",
		X"06",X"B7",X"11",X"04",X"00",X"ED",X"52",X"CD",X"C6",X"04",X"21",X"A1",X"80",X"35",X"20",X"E4",
		X"36",X"20",X"21",X"A5",X"80",X"34",X"18",X"DC",X"2A",X"A7",X"80",X"11",X"50",X"00",X"3A",X"A6",
		X"80",X"E6",X"01",X"20",X"1B",X"B7",X"ED",X"52",X"22",X"A7",X"80",X"CD",X"C6",X"04",X"21",X"A2",
		X"80",X"35",X"20",X"06",X"36",X"10",X"21",X"A6",X"80",X"34",X"21",X"A5",X"80",X"35",X"18",X"B4",
		X"19",X"18",X"E5",X"3E",X"FF",X"C9",X"CD",X"C7",X"06",X"3E",X"18",X"32",X"B0",X"80",X"21",X"00",
		X"01",X"22",X"B1",X"80",X"AF",X"32",X"B3",X"80",X"21",X"00",X"02",X"22",X"B4",X"80",X"16",X"06",
		X"1E",X"00",X"CD",X"4C",X"05",X"CD",X"80",X"05",X"06",X"03",X"CD",X"FE",X"05",X"C9",X"2A",X"B4",
		X"80",X"2B",X"7C",X"B5",X"28",X"4B",X"22",X"B4",X"80",X"3A",X"B3",X"80",X"FE",X"00",X"28",X"1B",
		X"2A",X"B1",X"80",X"2B",X"7C",X"B5",X"20",X"34",X"21",X"00",X"01",X"22",X"B1",X"80",X"16",X"06",
		X"1E",X"00",X"CD",X"4C",X"05",X"AF",X"32",X"B3",X"80",X"AF",X"C9",X"21",X"B0",X"80",X"35",X"20",
		X"F8",X"36",X"18",X"16",X"06",X"CD",X"35",X"06",X"1C",X"7B",X"FE",X"08",X"28",X"05",X"CD",X"4C",
		X"05",X"18",X"E6",X"CD",X"4C",X"05",X"21",X"B3",X"80",X"34",X"18",X"DD",X"22",X"B1",X"80",X"18",
		X"D8",X"3E",X"FF",X"C9",X"CD",X"BC",X"07",X"3E",X"01",X"32",X"C0",X"80",X"21",X"00",X"08",X"22",
		X"C3",X"80",X"AF",X"32",X"C5",X"80",X"21",X"00",X"02",X"22",X"C6",X"80",X"21",X"00",X"05",X"CD",
		X"C6",X"04",X"CD",X"0D",X"05",X"06",X"08",X"CD",X"FE",X"05",X"C9",X"2A",X"C6",X"80",X"2B",X"7C",
		X"B5",X"28",X"43",X"22",X"C6",X"80",X"21",X"C0",X"80",X"35",X"20",X"2C",X"36",X"01",X"CD",X"80",
		X"06",X"11",X"08",X"00",X"19",X"ED",X"5B",X"C3",X"80",X"7C",X"BA",X"20",X"18",X"7D",X"BB",X"20",
		X"14",X"3A",X"C5",X"80",X"B7",X"20",X"13",X"21",X"00",X"0B",X"22",X"C3",X"80",X"3E",X"FF",X"32",
		X"C5",X"80",X"21",X"00",X"05",X"CD",X"C6",X"04",X"AF",X"C9",X"21",X"00",X"08",X"22",X"C3",X"80",
		X"AF",X"32",X"C5",X"80",X"18",X"EC",X"3E",X"FF",X"C9",X"CD",X"48",X"07",X"3E",X"08",X"32",X"D0",
		X"80",X"3E",X"05",X"32",X"D1",X"80",X"3E",X"0C",X"32",X"D2",X"80",X"AF",X"32",X"D3",X"80",X"21",
		X"50",X"00",X"CD",X"C6",X"04",X"CD",X"0D",X"05",X"06",X"00",X"CD",X"FE",X"05",X"C9",X"3A",X"D3",
		X"80",X"FE",X"00",X"28",X"18",X"FE",X"01",X"28",X"26",X"FE",X"02",X"28",X"27",X"FE",X"03",X"28",
		X"33",X"21",X"D2",X"80",X"35",X"28",X"32",X"AF",X"32",X"D3",X"80",X"AF",X"C9",X"CD",X"4B",X"06",
		X"3C",X"FE",X"0A",X"20",X"04",X"21",X"D3",X"80",X"34",X"47",X"CD",X"FE",X"05",X"18",X"EC",X"CD",
		X"1C",X"14",X"18",X"E7",X"CD",X"4B",X"06",X"3D",X"20",X"04",X"21",X"D3",X"80",X"34",X"47",X"CD",
		X"FE",X"05",X"18",X"D7",X"CD",X"29",X"14",X"18",X"D2",X"3E",X"FF",X"C9",X"21",X"D0",X"80",X"35",
		X"C0",X"3E",X"08",X"77",X"21",X"D3",X"80",X"34",X"C9",X"21",X"D1",X"80",X"35",X"C0",X"3E",X"05",
		X"77",X"21",X"D3",X"80",X"34",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
